
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_LWC_1 is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_LWC_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_LWC_1.all;

entity CryptoCore_1_DW01_cmp6_0 is

   port( A, B : in std_logic_vector (31 downto 0);  TC : in std_logic;  LT, GT,
         EQ, LE, GE, NE : out std_logic);

end CryptoCore_1_DW01_cmp6_0;

architecture SYN_rpl of CryptoCore_1_DW01_cmp6_0 is

   component NOR4X0
      port( IN1, IN2, IN3, IN4 : in std_logic;  QN : out std_logic);
   end component;
   
   component NOR2X0
      port( IN1, IN2 : in std_logic;  QN : out std_logic);
   end component;
   
   component OA22X1
      port( IN1, IN2, IN3, IN4 : in std_logic;  Q : out std_logic);
   end component;
   
   component AND2X1
      port( IN1, IN2 : in std_logic;  Q : out std_logic);
   end component;
   
   component XNOR2X1
      port( IN1, IN2 : in std_logic;  Q : out std_logic);
   end component;
   
   component NAND4X0
      port( IN1, IN2, IN3, IN4 : in std_logic;  QN : out std_logic);
   end component;
   
   component INVX0
      port( INP : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2X2
      port( IN1, IN2 : in std_logic;  Q : out std_logic);
   end component;
   
   component XNOR2X2
      port( IN1, IN2 : in std_logic;  Q : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49 : std_logic;

begin
   
   U1 : INVX0 port map( INP => A(3), ZN => n1);
   U2 : INVX0 port map( INP => A(2), ZN => n2);
   U3 : NOR4X0 port map( IN1 => n40, IN2 => n41, IN3 => n42, IN4 => n43, QN => 
                           n7);
   U4 : XNOR2X2 port map( IN1 => B(14), IN2 => A(14), Q => n33);
   U5 : XNOR2X2 port map( IN1 => B(15), IN2 => A(15), Q => n32);
   U6 : XNOR2X1 port map( IN1 => B(3), IN2 => n1, Q => n43);
   U7 : XNOR2X1 port map( IN1 => B(2), IN2 => n2, Q => n42);
   U8 : XNOR2X2 port map( IN1 => B(23), IN2 => A(23), Q => n22);
   U9 : XNOR2X2 port map( IN1 => B(26), IN2 => A(26), Q => n19);
   U10 : XNOR2X2 port map( IN1 => B(13), IN2 => A(13), Q => n34);
   U11 : XNOR2X2 port map( IN1 => B(20), IN2 => A(20), Q => n25);
   U12 : XNOR2X2 port map( IN1 => B(30), IN2 => A(30), Q => n15);
   U13 : INVX0 port map( INP => A(1), ZN => n4);
   U14 : INVX0 port map( INP => A(0), ZN => n5);
   U15 : XNOR2X2 port map( IN1 => B(19), IN2 => A(19), Q => n26);
   U16 : XNOR2X2 port map( IN1 => B(9), IN2 => A(9), Q => n38);
   U17 : XNOR2X2 port map( IN1 => B(18), IN2 => A(18), Q => n27);
   U18 : XNOR2X2 port map( IN1 => B(16), IN2 => A(16), Q => n29);
   U19 : XNOR2X2 port map( IN1 => B(21), IN2 => A(21), Q => n24);
   U20 : XNOR2X2 port map( IN1 => B(27), IN2 => A(27), Q => n18);
   U21 : XNOR2X2 port map( IN1 => B(24), IN2 => A(24), Q => n21);
   U22 : XNOR2X2 port map( IN1 => B(31), IN2 => A(31), Q => n14);
   U23 : XOR2X2 port map( IN1 => B(7), IN2 => A(7), Q => n49);
   U24 : XNOR2X2 port map( IN1 => B(29), IN2 => A(29), Q => n16);
   U25 : XNOR2X2 port map( IN1 => B(25), IN2 => A(25), Q => n20);
   U26 : XNOR2X2 port map( IN1 => B(28), IN2 => A(28), Q => n17);
   U27 : XOR2X2 port map( IN1 => B(4), IN2 => A(4), Q => n46);
   U28 : XOR2X2 port map( IN1 => B(5), IN2 => A(5), Q => n47);
   U29 : XOR2X2 port map( IN1 => B(6), IN2 => A(6), Q => n48);
   U30 : INVX0 port map( INP => B(1), ZN => n3);
   U31 : NAND4X0 port map( IN1 => n9, IN2 => n7, IN3 => n8, IN4 => n6, QN => NE
                           );
   U32 : NOR4X0 port map( IN1 => n10, IN2 => n11, IN3 => n12, IN4 => n13, QN =>
                           n9);
   U33 : NAND4X0 port map( IN1 => n14, IN2 => n15, IN3 => n16, IN4 => n17, QN 
                           => n13);
   U34 : NAND4X0 port map( IN1 => n18, IN2 => n19, IN3 => n20, IN4 => n21, QN 
                           => n12);
   U35 : NAND4X0 port map( IN1 => n22, IN2 => n23, IN3 => n24, IN4 => n25, QN 
                           => n11);
   U36 : XNOR2X1 port map( IN1 => B(22), IN2 => A(22), Q => n23);
   U37 : NAND4X0 port map( IN1 => n26, IN2 => n27, IN3 => n28, IN4 => n29, QN 
                           => n10);
   U38 : XNOR2X1 port map( IN1 => B(17), IN2 => A(17), Q => n28);
   U39 : NOR2X0 port map( IN1 => n31, IN2 => n30, QN => n8);
   U40 : NAND4X0 port map( IN1 => n32, IN2 => n33, IN3 => n34, IN4 => n35, QN 
                           => n31);
   U41 : XNOR2X1 port map( IN1 => B(12), IN2 => A(12), Q => n35);
   U42 : NAND4X0 port map( IN1 => n36, IN2 => n37, IN3 => n38, IN4 => n39, QN 
                           => n30);
   U43 : XNOR2X1 port map( IN1 => B(8), IN2 => A(8), Q => n39);
   U44 : XNOR2X1 port map( IN1 => B(10), IN2 => A(10), Q => n37);
   U45 : XNOR2X1 port map( IN1 => B(11), IN2 => A(11), Q => n36);
   U46 : OA22X1 port map( IN1 => B(1), IN2 => n44, IN3 => n44, IN4 => n4, Q => 
                           n41);
   U47 : AND2X1 port map( IN1 => B(0), IN2 => n5, Q => n44);
   U48 : OA22X1 port map( IN1 => n45, IN2 => n3, IN3 => A(1), IN4 => n45, Q => 
                           n40);
   U49 : NOR2X0 port map( IN1 => n5, IN2 => B(0), QN => n45);
   U50 : NOR4X0 port map( IN1 => n46, IN2 => n47, IN3 => n48, IN4 => n49, QN =>
                           n6);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_LWC_1.all;

entity counter_num_bits4_1_1 is

   port( clk, load, enable : in std_logic;  start_value : in std_logic_vector 
         (3 downto 0);  q : out std_logic_vector (3 downto 0));

end counter_num_bits4_1_1;

architecture SYN_Behavioral of counter_num_bits4_1_1 is

   component NOR2X0
      port( IN1, IN2 : in std_logic;  QN : out std_logic);
   end component;
   
   component INVX0
      port( INP : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4X0
      port( IN1, IN2, IN3, IN4 : in std_logic;  QN : out std_logic);
   end component;
   
   component AO222X1
      port( IN1, IN2, IN3, IN4, IN5, IN6 : in std_logic;  Q : out std_logic);
   end component;
   
   component NAND3X0
      port( IN1, IN2, IN3 : in std_logic;  QN : out std_logic);
   end component;
   
   component OAI21X1
      port( IN1, IN2, IN3 : in std_logic;  QN : out std_logic);
   end component;
   
   component AO21X1
      port( IN1, IN2, IN3 : in std_logic;  Q : out std_logic);
   end component;
   
   component AO221X1
      port( IN1, IN2, IN3, IN4, IN5 : in std_logic;  Q : out std_logic);
   end component;
   
   component DFFX1
      port( D, CLK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal q_3_port, q_2_port, q_1_port, q_0_port, n3, n4, n5, n18, n19, n20, 
      n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n_1006, n_1007 : 
      std_logic;

begin
   q <= ( q_3_port, q_2_port, q_1_port, q_0_port );
   
   count_reg_0_inst : DFFX1 port map( D => n18, CLK => clk, Q => q_0_port, QN 
                           => n_1006);
   count_reg_1_inst : DFFX1 port map( D => n19, CLK => clk, Q => q_1_port, QN 
                           => n30);
   count_reg_2_inst : DFFX1 port map( D => n20, CLK => clk, Q => q_2_port, QN 
                           => n31);
   count_reg_3_inst : DFFX1 port map( D => n21, CLK => clk, Q => q_3_port, QN 
                           => n_1007);
   U10 : AO221X1 port map( IN1 => q_3_port, IN2 => n29, IN3 => start_value(3), 
                           IN4 => load, IN5 => n28, Q => n21);
   U11 : AO21X1 port map( IN1 => n4, IN2 => n31, IN3 => n26, Q => n29);
   U12 : AO222X1 port map( IN1 => start_value(2), IN2 => load, IN3 => n25, IN4 
                           => q_1_port, IN5 => q_2_port, IN6 => n26, Q => n20);
   U13 : AO21X1 port map( IN1 => n4, IN2 => n30, IN3 => n24, Q => n26);
   U14 : AO222X1 port map( IN1 => n3, IN2 => n30, IN3 => start_value(1), IN4 =>
                           load, IN5 => q_1_port, IN6 => n24, Q => n19);
   U15 : OAI21X1 port map( IN1 => load, IN2 => q_0_port, IN3 => n5, QN => n24);
   U16 : NAND3X0 port map( IN1 => n5, IN2 => n4, IN3 => q_0_port, QN => n27);
   U17 : AO222X1 port map( IN1 => start_value(0), IN2 => load, IN3 => n23, IN4 
                           => n5, IN5 => n22, IN6 => q_0_port, Q => n18);
   U3 : INVX0 port map( INP => n22, ZN => n5);
   U4 : INVX0 port map( INP => load, ZN => n4);
   U5 : NOR2X0 port map( IN1 => enable, IN2 => load, QN => n22);
   U6 : NOR4X0 port map( IN1 => q_3_port, IN2 => n27, IN3 => n30, IN4 => n31, 
                           QN => n28);
   U7 : INVX0 port map( INP => n27, ZN => n3);
   U8 : NOR2X0 port map( IN1 => q_2_port, IN2 => n27, QN => n25);
   U9 : NOR2X0 port map( IN1 => q_0_port, IN2 => load, QN => n23);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_LWC_1.all;

entity StepDownCountLd_N16_step4_1_1 is

   port( clk, len, ena : in std_logic;  load : in std_logic_vector (15 downto 
         0);  count : out std_logic_vector (15 downto 0));

end StepDownCountLd_N16_step4_1_1;

architecture SYN_StepDownCountLd of StepDownCountLd_N16_step4_1_1 is

   component XNOR2X1
      port( IN1, IN2 : in std_logic;  Q : out std_logic);
   end component;
   
   component OR2X1
      port( IN1, IN2 : in std_logic;  Q : out std_logic);
   end component;
   
   component NOR2X0
      port( IN1, IN2 : in std_logic;  QN : out std_logic);
   end component;
   
   component NBUFFX2
      port( INP : in std_logic;  Z : out std_logic);
   end component;
   
   component AO222X1
      port( IN1, IN2, IN3, IN4, IN5, IN6 : in std_logic;  Q : out std_logic);
   end component;
   
   component DFFX1
      port( D, CLK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal count_15_port, count_14_port, count_13_port, count_12_port, 
      count_11_port, count_10_port, count_9_port, count_8_port, count_7_port, 
      count_6_port, count_5_port, count_4_port, count_3_port, count_2_port, N4,
      N5, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18, N19, 
      sub_55_carry_4_port, sub_55_carry_5_port, sub_55_carry_6_port, 
      sub_55_carry_7_port, sub_55_carry_8_port, sub_55_carry_9_port, 
      sub_55_carry_10_port, sub_55_carry_11_port, sub_55_carry_12_port, 
      sub_55_carry_13_port, sub_55_carry_14_port, sub_55_carry_15_port, n1, n2,
      n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35
      , n36, n37, n38, n39, n_1008, n_1009, n_1010, n_1011, n_1012, n_1013, 
      n_1014, n_1015, n_1016, n_1017, n_1018, n_1019, n_1020, n_1021, n_1022 : 
      std_logic;

begin
   count <= ( count_15_port, count_14_port, count_13_port, count_12_port, 
      count_11_port, count_10_port, count_9_port, count_8_port, count_7_port, 
      count_6_port, count_5_port, count_4_port, count_3_port, count_2_port, N5,
      N4 );
   
   qtemp_reg_0_inst : DFFX1 port map( D => n22, CLK => clk, Q => N4, QN => 
                           n_1008);
   qtemp_reg_1_inst : DFFX1 port map( D => n23, CLK => clk, Q => N5, QN => 
                           n_1009);
   qtemp_reg_2_inst : DFFX1 port map( D => n24, CLK => clk, Q => count_2_port, 
                           QN => n1);
   qtemp_reg_3_inst : DFFX1 port map( D => n25, CLK => clk, Q => count_3_port, 
                           QN => n_1010);
   qtemp_reg_4_inst : DFFX1 port map( D => n26, CLK => clk, Q => count_4_port, 
                           QN => n_1011);
   qtemp_reg_5_inst : DFFX1 port map( D => n27, CLK => clk, Q => count_5_port, 
                           QN => n_1012);
   qtemp_reg_6_inst : DFFX1 port map( D => n28, CLK => clk, Q => count_6_port, 
                           QN => n_1013);
   qtemp_reg_7_inst : DFFX1 port map( D => n29, CLK => clk, Q => count_7_port, 
                           QN => n_1014);
   qtemp_reg_8_inst : DFFX1 port map( D => n30, CLK => clk, Q => count_8_port, 
                           QN => n_1015);
   qtemp_reg_9_inst : DFFX1 port map( D => n31, CLK => clk, Q => count_9_port, 
                           QN => n_1016);
   qtemp_reg_10_inst : DFFX1 port map( D => n32, CLK => clk, Q => count_10_port
                           , QN => n_1017);
   qtemp_reg_11_inst : DFFX1 port map( D => n33, CLK => clk, Q => count_11_port
                           , QN => n_1018);
   qtemp_reg_12_inst : DFFX1 port map( D => n34, CLK => clk, Q => count_12_port
                           , QN => n_1019);
   qtemp_reg_13_inst : DFFX1 port map( D => n35, CLK => clk, Q => count_13_port
                           , QN => n_1020);
   qtemp_reg_14_inst : DFFX1 port map( D => n36, CLK => clk, Q => count_14_port
                           , QN => n_1021);
   qtemp_reg_15_inst : DFFX1 port map( D => n37, CLK => clk, Q => count_15_port
                           , QN => n_1022);
   U6 : AO222X1 port map( IN1 => load(15), IN2 => n21, IN3 => N19, IN4 => n39, 
                           IN5 => count_15_port, IN6 => n38, Q => n37);
   U7 : AO222X1 port map( IN1 => load(14), IN2 => n21, IN3 => N18, IN4 => n39, 
                           IN5 => count_14_port, IN6 => n38, Q => n36);
   U8 : AO222X1 port map( IN1 => load(13), IN2 => n21, IN3 => N17, IN4 => n39, 
                           IN5 => count_13_port, IN6 => n38, Q => n35);
   U9 : AO222X1 port map( IN1 => load(12), IN2 => n21, IN3 => N16, IN4 => n39, 
                           IN5 => count_12_port, IN6 => n38, Q => n34);
   U10 : AO222X1 port map( IN1 => load(11), IN2 => n21, IN3 => N15, IN4 => n39,
                           IN5 => count_11_port, IN6 => n38, Q => n33);
   U11 : AO222X1 port map( IN1 => load(10), IN2 => n21, IN3 => N14, IN4 => n39,
                           IN5 => count_10_port, IN6 => n38, Q => n32);
   U12 : AO222X1 port map( IN1 => load(9), IN2 => n21, IN3 => N13, IN4 => n39, 
                           IN5 => count_9_port, IN6 => n38, Q => n31);
   U13 : AO222X1 port map( IN1 => load(8), IN2 => n21, IN3 => N12, IN4 => n39, 
                           IN5 => count_8_port, IN6 => n38, Q => n30);
   U14 : AO222X1 port map( IN1 => load(7), IN2 => n21, IN3 => N11, IN4 => n39, 
                           IN5 => count_7_port, IN6 => n38, Q => n29);
   U15 : AO222X1 port map( IN1 => load(6), IN2 => n21, IN3 => N10, IN4 => n39, 
                           IN5 => count_6_port, IN6 => n38, Q => n28);
   U16 : AO222X1 port map( IN1 => load(5), IN2 => n21, IN3 => N9, IN4 => n39, 
                           IN5 => count_5_port, IN6 => n38, Q => n27);
   U17 : AO222X1 port map( IN1 => load(4), IN2 => n21, IN3 => N8, IN4 => n39, 
                           IN5 => count_4_port, IN6 => n38, Q => n26);
   U18 : AO222X1 port map( IN1 => load(3), IN2 => n21, IN3 => N7, IN4 => n39, 
                           IN5 => count_3_port, IN6 => n38, Q => n25);
   U19 : AO222X1 port map( IN1 => load(2), IN2 => n21, IN3 => n1, IN4 => n39, 
                           IN5 => count_2_port, IN6 => n38, Q => n24);
   U20 : AO222X1 port map( IN1 => load(1), IN2 => n21, IN3 => N5, IN4 => n39, 
                           IN5 => N5, IN6 => n38, Q => n23);
   U21 : AO222X1 port map( IN1 => load(0), IN2 => n21, IN3 => N4, IN4 => n39, 
                           IN5 => N4, IN6 => n38, Q => n22);
   U3 : NOR2X0 port map( IN1 => n38, IN2 => n2, QN => n39);
   U4 : NBUFFX2 port map( INP => len, Z => n21);
   U5 : NBUFFX2 port map( INP => len, Z => n2);
   U22 : NOR2X0 port map( IN1 => ena, IN2 => n2, QN => n38);
   U23 : XNOR2X1 port map( IN1 => sub_55_carry_15_port, IN2 => count_15_port, Q
                           => N19);
   U24 : OR2X1 port map( IN1 => sub_55_carry_14_port, IN2 => count_14_port, Q 
                           => sub_55_carry_15_port);
   U25 : XNOR2X1 port map( IN1 => count_14_port, IN2 => sub_55_carry_14_port, Q
                           => N18);
   U26 : OR2X1 port map( IN1 => sub_55_carry_13_port, IN2 => count_13_port, Q 
                           => sub_55_carry_14_port);
   U27 : XNOR2X1 port map( IN1 => count_13_port, IN2 => sub_55_carry_13_port, Q
                           => N17);
   U28 : OR2X1 port map( IN1 => sub_55_carry_12_port, IN2 => count_12_port, Q 
                           => sub_55_carry_13_port);
   U29 : XNOR2X1 port map( IN1 => count_12_port, IN2 => sub_55_carry_12_port, Q
                           => N16);
   U30 : OR2X1 port map( IN1 => sub_55_carry_11_port, IN2 => count_11_port, Q 
                           => sub_55_carry_12_port);
   U31 : XNOR2X1 port map( IN1 => count_11_port, IN2 => sub_55_carry_11_port, Q
                           => N15);
   U32 : OR2X1 port map( IN1 => sub_55_carry_10_port, IN2 => count_10_port, Q 
                           => sub_55_carry_11_port);
   U33 : XNOR2X1 port map( IN1 => count_10_port, IN2 => sub_55_carry_10_port, Q
                           => N14);
   U34 : OR2X1 port map( IN1 => sub_55_carry_9_port, IN2 => count_9_port, Q => 
                           sub_55_carry_10_port);
   U35 : XNOR2X1 port map( IN1 => count_9_port, IN2 => sub_55_carry_9_port, Q 
                           => N13);
   U36 : OR2X1 port map( IN1 => sub_55_carry_8_port, IN2 => count_8_port, Q => 
                           sub_55_carry_9_port);
   U37 : XNOR2X1 port map( IN1 => count_8_port, IN2 => sub_55_carry_8_port, Q 
                           => N12);
   U38 : OR2X1 port map( IN1 => sub_55_carry_7_port, IN2 => count_7_port, Q => 
                           sub_55_carry_8_port);
   U39 : XNOR2X1 port map( IN1 => count_7_port, IN2 => sub_55_carry_7_port, Q 
                           => N11);
   U40 : OR2X1 port map( IN1 => sub_55_carry_6_port, IN2 => count_6_port, Q => 
                           sub_55_carry_7_port);
   U41 : XNOR2X1 port map( IN1 => count_6_port, IN2 => sub_55_carry_6_port, Q 
                           => N10);
   U42 : OR2X1 port map( IN1 => sub_55_carry_5_port, IN2 => count_5_port, Q => 
                           sub_55_carry_6_port);
   U43 : XNOR2X1 port map( IN1 => count_5_port, IN2 => sub_55_carry_5_port, Q 
                           => N9);
   U44 : OR2X1 port map( IN1 => sub_55_carry_4_port, IN2 => count_4_port, Q => 
                           sub_55_carry_5_port);
   U45 : XNOR2X1 port map( IN1 => count_4_port, IN2 => sub_55_carry_4_port, Q 
                           => N8);
   U46 : OR2X1 port map( IN1 => count_2_port, IN2 => count_3_port, Q => 
                           sub_55_carry_4_port);
   U47 : XNOR2X1 port map( IN1 => count_3_port, IN2 => count_2_port, Q => N7);

end SYN_StepDownCountLd;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_LWC_1.all;

entity DATA_SIPO_1 is

   port( clk, rst, end_of_input : in std_logic;  data_p : out std_logic_vector 
         (31 downto 0);  data_valid_p : out std_logic;  data_ready_p : in 
         std_logic;  data_s : in std_logic_vector (31 downto 0);  data_valid_s 
         : in std_logic;  data_ready_s : out std_logic);

end DATA_SIPO_1;

architecture SYN_behavioral of DATA_SIPO_1 is

begin
   data_p <= ( data_s(31), data_s(30), data_s(29), data_s(28), data_s(27), 
      data_s(26), data_s(25), data_s(24), data_s(23), data_s(22), data_s(21), 
      data_s(20), data_s(19), data_s(18), data_s(17), data_s(16), data_s(15), 
      data_s(14), data_s(13), data_s(12), data_s(11), data_s(10), data_s(9), 
      data_s(8), data_s(7), data_s(6), data_s(5), data_s(4), data_s(3), 
      data_s(2), data_s(1), data_s(0) );
   data_valid_p <= data_valid_s;
   data_ready_s <= data_ready_p;

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_LWC_1.all;

entity cyclist_ops_RAM_LEN128_DATA_LEN32_1 is

   port( cyc_state_update_sel, xor_sel, cycd_sel : in std_logic_vector (1 
         downto 0);  extract_sel, addr_sel2 : in std_logic;  ramoutd1 : in 
         std_logic_vector (127 downto 0);  key, bdi_data : in std_logic_vector 
         (31 downto 0);  cu_cd : in std_logic_vector (7 downto 0);  dcount_in :
         in std_logic_vector (1 downto 0);  cyc_state_update : out 
         std_logic_vector (127 downto 0);  bdo_out : out std_logic_vector (31 
         downto 0));

end cyclist_ops_RAM_LEN128_DATA_LEN32_1;

architecture SYN_Behavioral of cyclist_ops_RAM_LEN128_DATA_LEN32_1 is

   component NOR2X0
      port( IN1, IN2 : in std_logic;  QN : out std_logic);
   end component;
   
   component NAND2X0
      port( IN1, IN2 : in std_logic;  QN : out std_logic);
   end component;
   
   component INVX0
      port( INP : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2X1
      port( IN1, IN2 : in std_logic;  Q : out std_logic);
   end component;
   
   component NBUFFX2
      port( INP : in std_logic;  Z : out std_logic);
   end component;
   
   component AO22X1
      port( IN1, IN2, IN3, IN4 : in std_logic;  Q : out std_logic);
   end component;
   
   component XOR2X1
      port( IN1, IN2 : in std_logic;  Q : out std_logic);
   end component;
   
   component OR2X1
      port( IN1, IN2 : in std_logic;  Q : out std_logic);
   end component;
   
   component NAND2X1
      port( IN1, IN2 : in std_logic;  QN : out std_logic);
   end component;
   
   component AO22X2
      port( IN1, IN2, IN3, IN4 : in std_logic;  Q : out std_logic);
   end component;
   
   component DELLN2X2
      port( INP : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3X0
      port( IN1, IN2, IN3 : in std_logic;  QN : out std_logic);
   end component;
   
   component IBUFFX16
      port( INP : in std_logic;  ZN : out std_logic);
   end component;
   
   component AO221X1
      port( IN1, IN2, IN3, IN4, IN5 : in std_logic;  Q : out std_logic);
   end component;
   
   component MUX41X1
      port( IN1, IN3, IN2, IN4, S0, S1 : in std_logic;  Q : out std_logic);
   end component;
   
   component AO222X1
      port( IN1, IN2, IN3, IN4, IN5, IN6 : in std_logic;  Q : out std_logic);
   end component;
   
   component DELLN1X2
      port( INP : in std_logic;  Z : out std_logic);
   end component;
   
   component AO221X2
      port( IN1, IN2, IN3, IN4, IN5 : in std_logic;  Q : out std_logic);
   end component;
   
   component NOR2X4
      port( IN1, IN2 : in std_logic;  QN : out std_logic);
   end component;
   
   component NOR2X1
      port( IN1, IN2 : in std_logic;  QN : out std_logic);
   end component;
   
   component NAND2X2
      port( IN1, IN2 : in std_logic;  QN : out std_logic);
   end component;
   
   component MUX41X2
      port( IN1, IN3, IN2, IN4, S0, S1 : in std_logic;  Q : out std_logic);
   end component;
   
   component NBUFFX32
      port( INP : in std_logic;  Z : out std_logic);
   end component;
   
   component INVX4
      port( INP : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2X4
      port( IN1, IN2 : in std_logic;  QN : out std_logic);
   end component;
   
   component AO21X1
      port( IN1, IN2, IN3 : in std_logic;  Q : out std_logic);
   end component;
   
   component XNOR2X1
      port( IN1, IN2 : in std_logic;  Q : out std_logic);
   end component;
   
   component OA21X1
      port( IN1, IN2, IN3 : in std_logic;  Q : out std_logic);
   end component;
   
   signal n18, n19, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
      n33, n35, n36, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49
      , n50, n51, n52, n53, n54, n56, n57, n58, n59, n60, n61, n62, n63, n64, 
      n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79
      , n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, 
      n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, 
      n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, 
      n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, 
      n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, 
      n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n155, 
      n156, n157, n158, n159, n160, n161, n162, n164, n165, n166, n168, n169, 
      n171, n172, n174, n175, n177, n178, n179, n180, n181, n182, n183, n184, 
      n186, n187, n188, n189, n191, n192, n193, n194, n195, n196, n197, n198, 
      n199, n201, n202, n204, n206, n208, n209, n211, n213, n215, n217, n218, 
      n221, n223, n225, n227, n229, n231, n232, n233, n234, n1, n2, n3, n4, n5,
      n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n20, n34, n37, 
      n55, n154, n163, n167, n170, n173, n176, n185, n190, n200, n203, n205, 
      n207, n210, n212, n214, n216, n219, n220, n222, n224, n226, n228, n230, 
      n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, 
      n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, 
      n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, 
      n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, 
      n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, 
      n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, 
      n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, 
      n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, 
      n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, 
      n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, 
      n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, 
      n367, n368, n369, n370, n371, n372, n373 : std_logic;

begin
   
   U46 : AO22X1 port map( IN1 => n314, IN2 => n21, IN3 => n325, IN4 => n347, Q 
                           => cyc_state_update(99));
   U51 : AO22X1 port map( IN1 => n306, IN2 => n28, IN3 => ramoutd1(94), IN4 => 
                           n344, Q => cyc_state_update(94));
   U52 : AO22X1 port map( IN1 => n306, IN2 => n247, IN3 => n280, IN4 => n344, Q
                           => cyc_state_update(93));
   U54 : AO22X1 port map( IN1 => n307, IN2 => n31, IN3 => n270, IN4 => n344, Q 
                           => cyc_state_update(91));
   U61 : AO22X1 port map( IN1 => n239, IN2 => n309, IN3 => ramoutd1(85), IN4 =>
                           n344, Q => cyc_state_update(85));
   U62 : AO22X1 port map( IN1 => n309, IN2 => n39, IN3 => ramoutd1(84), IN4 => 
                           n344, Q => cyc_state_update(84));
   U66 : AO22X1 port map( IN1 => n308, IN2 => n43, IN3 => ramoutd1(80), IN4 => 
                           n345, Q => cyc_state_update(80));
   U67 : AO22X1 port map( IN1 => n302, IN2 => n44, IN3 => ramoutd1(7), IN4 => 
                           n351, Q => cyc_state_update(7));
   U69 : AO22X1 port map( IN1 => n308, IN2 => n46, IN3 => n55, IN4 => n345, Q 
                           => cyc_state_update(78));
   U73 : AO22X1 port map( IN1 => n308, IN2 => n190, IN3 => ramoutd1(74), IN4 =>
                           n345, Q => cyc_state_update(74));
   U76 : AO22X1 port map( IN1 => n307, IN2 => n44, IN3 => n261, IN4 => n346, Q 
                           => cyc_state_update(71));
   U92 : AO22X1 port map( IN1 => n311, IN2 => n15, IN3 => ramoutd1(57), IN4 => 
                           n340, Q => cyc_state_update(57));
   U100 : AO22X1 port map( IN1 => n303, IN2 => n53, IN3 => n319, IN4 => n351, Q
                           => cyc_state_update(4));
   U104 : AO22X1 port map( IN1 => n312, IN2 => n241, IN3 => ramoutd1(46), IN4 
                           => n341, Q => cyc_state_update(46));
   U112 : AO22X1 port map( IN1 => n312, IN2 => n44, IN3 => ramoutd1(39), IN4 =>
                           n342, Q => cyc_state_update(39));
   U117 : AO222X1 port map( IN1 => key(3), IN2 => n339, IN3 => bdi_data(3), IN4
                           => n360, IN5 => n334, IN6 => n59, Q => n21);
   U119 : AO22X1 port map( IN1 => n313, IN2 => n24, IN3 => ramoutd1(33), IN4 =>
                           n342, Q => cyc_state_update(33));
   U124 : AO222X1 port map( IN1 => key(2), IN2 => n338, IN3 => bdi_data(2), IN4
                           => n360, IN5 => n334, IN6 => n62, Q => n23);
   U136 : AO222X1 port map( IN1 => key(1), IN2 => n338, IN3 => bdi_data(1), IN4
                           => n360, IN5 => n334, IN6 => n63, Q => n24);
   U146 : AO221X1 port map( IN1 => key(31), IN2 => n338, IN3 => n64, IN4 => 
                           n334, IN5 => n65, Q => n26);
   U149 : AO221X1 port map( IN1 => key(30), IN2 => n338, IN3 => n69, IN4 => 
                           n336, IN5 => n70, Q => n28);
   U152 : AO221X1 port map( IN1 => key(29), IN2 => n338, IN3 => n72, IN4 => 
                           n336, IN5 => n73, Q => n29);
   U155 : AO221X1 port map( IN1 => key(28), IN2 => n338, IN3 => n75, IN4 => 
                           n336, IN5 => n76, Q => n30);
   U159 : AO22X1 port map( IN1 => bdi_data(27), IN2 => n66, IN3 => n67, IN4 => 
                           n269, Q => n79);
   U161 : AO221X1 port map( IN1 => key(26), IN2 => n337, IN3 => n81, IN4 => 
                           n335, IN5 => n82, Q => n32);
   U166 : OA21X1 port map( IN1 => n363, IN2 => n87, IN3 => n360, Q => n67);
   U167 : AND2X1 port map( IN1 => n88, IN2 => n360, Q => n66);
   U169 : AO222X1 port map( IN1 => key(24), IN2 => n338, IN3 => n360, IN4 => 
                           n89, IN5 => n334, IN6 => n90, Q => n35);
   U170 : AO222X1 port map( IN1 => bdi_data(24), IN2 => n88, IN3 => n363, IN4 
                           => n264, IN5 => n87, IN6 => n367, Q => n89);
   U173 : AO221X1 port map( IN1 => key(23), IN2 => n338, IN3 => n93, IN4 => 
                           n335, IN5 => n94, Q => n36);
   U174 : AO22X1 port map( IN1 => bdi_data(23), IN2 => n95, IN3 => n96, IN4 => 
                           n97, Q => n94);
   U178 : AO22X1 port map( IN1 => n316, IN2 => n239, IN3 => n318, IN4 => n348, 
                           Q => cyc_state_update(117));
   U179 : AO221X1 port map( IN1 => key(21), IN2 => n337, IN3 => n101, IN4 => 
                           n335, IN5 => n102, Q => n38);
   U181 : AO22X1 port map( IN1 => n316, IN2 => n39, IN3 => ramoutd1(116), IN4 
                           => n348, Q => cyc_state_update(116));
   U182 : AO221X1 port map( IN1 => key(20), IN2 => n337, IN3 => n104, IN4 => 
                           n335, IN5 => n105, Q => n39);
   U184 : AO22X1 port map( IN1 => n40, IN2 => n316, IN3 => n262, IN4 => n348, Q
                           => cyc_state_update(115));
   U185 : AO221X1 port map( IN1 => key(19), IN2 => n337, IN3 => n107, IN4 => 
                           n335, IN5 => n108, Q => n40);
   U188 : AO221X1 port map( IN1 => key(18), IN2 => n337, IN3 => n110, IN4 => 
                           n335, IN5 => n111, Q => n41);
   U191 : AO221X1 port map( IN1 => key(17), IN2 => n337, IN3 => n113, IN4 => 
                           n335, IN5 => n114, Q => n42);
   U193 : AO22X1 port map( IN1 => n316, IN2 => n43, IN3 => ramoutd1(112), IN4 
                           => n348, Q => cyc_state_update(112));
   U194 : AO222X1 port map( IN1 => key(16), IN2 => n338, IN3 => n360, IN4 => 
                           n119, IN5 => n334, IN6 => n120, Q => n43);
   U195 : AO222X1 port map( IN1 => n366, IN2 => n117, IN3 => bdi_data(16), IN4 
                           => n362, IN5 => n364, IN6 => n255, Q => n119);
   U197 : AO221X1 port map( IN1 => key(15), IN2 => n337, IN3 => n335, IN4 => 
                           n122, IN5 => n123, Q => n45);
   U198 : AO22X1 port map( IN1 => n124, IN2 => n125, IN3 => bdi_data(15), IN4 
                           => n126, Q => n123);
   U199 : AO22X1 port map( IN1 => n241, IN2 => n315, IN3 => n250, IN4 => n348, 
                           Q => cyc_state_update(110));
   U201 : AO22X1 port map( IN1 => n124, IN2 => n260, IN3 => bdi_data(14), IN4 
                           => n126, Q => n128);
   U204 : AO221X1 port map( IN1 => key(13), IN2 => n337, IN3 => n130, IN4 => 
                           n335, IN5 => n131, Q => n47);
   U205 : AO22X1 port map( IN1 => n124, IN2 => n185, IN3 => bdi_data(13), IN4 
                           => n126, Q => n131);
   U207 : AO221X1 port map( IN1 => key(12), IN2 => n337, IN3 => n133, IN4 => 
                           n335, IN5 => n134, Q => n48);
   U208 : AO22X1 port map( IN1 => n124, IN2 => n238, IN3 => bdi_data(12), IN4 
                           => n126, Q => n134);
   U210 : AO221X1 port map( IN1 => key(11), IN2 => n337, IN3 => n136, IN4 => 
                           n335, IN5 => n137, Q => n49);
   U211 : AO22X1 port map( IN1 => n124, IN2 => n220, IN3 => bdi_data(11), IN4 
                           => n126, Q => n137);
   U213 : AO221X1 port map( IN1 => key(10), IN2 => n337, IN3 => n335, IN4 => 
                           n139, IN5 => n140, Q => n50);
   U214 : AO22X1 port map( IN1 => n124, IN2 => n141, IN3 => bdi_data(10), IN4 
                           => n126, Q => n140);
   U216 : AO221X1 port map( IN1 => key(9), IN2 => n337, IN3 => n142, IN4 => 
                           n334, IN5 => n143, Q => n18);
   U217 : AO22X1 port map( IN1 => n124, IN2 => n13, IN3 => bdi_data(9), IN4 => 
                           n126, Q => n143);
   U218 : AO22X1 port map( IN1 => n246, IN2 => n317, IN3 => n4, IN4 => n349, Q 
                           => cyc_state_update(104));
   U219 : AO221X1 port map( IN1 => n334, IN2 => n145, IN3 => 
                           cyc_state_update_sel(1), IN4 => n361, IN5 => n146, Q
                           => n33);
   U220 : AO222X1 port map( IN1 => n368, IN2 => n124, IN3 => bdi_data(8), IN4 
                           => n126, IN5 => key(8), IN6 => n337, Q => n146);
   U221 : OA21X1 port map( IN1 => n362, IN2 => n117, IN3 => n360, Q => n126);
   U222 : AO22X1 port map( IN1 => n44, IN2 => n317, IN3 => n326, IN4 => n349, Q
                           => cyc_state_update(103));
   U223 : AO222X1 port map( IN1 => key(7), IN2 => n338, IN3 => bdi_data(7), IN4
                           => n360, IN5 => n334, IN6 => n148, Q => n44);
   U225 : AO222X1 port map( IN1 => key(6), IN2 => n339, IN3 => bdi_data(6), IN4
                           => n360, IN5 => n334, IN6 => n149, Q => n51);
   U227 : AO222X1 port map( IN1 => key(5), IN2 => n339, IN3 => bdi_data(5), IN4
                           => n360, IN5 => n334, IN6 => n150, Q => n52);
   U229 : AO222X1 port map( IN1 => key(4), IN2 => n339, IN3 => bdi_data(4), IN4
                           => n360, IN5 => n334, IN6 => n152, Q => n53);
   U231 : AO222X1 port map( IN1 => key(0), IN2 => n338, IN3 => bdi_data(0), IN4
                           => n360, IN5 => n334, IN6 => n153, Q => n25);
   U232 : AO22X1 port map( IN1 => n13, IN2 => n358, IN3 => n354, IN4 => n142, Q
                           => bdo_out(9));
   U237 : AO22X1 port map( IN1 => n263, IN2 => n358, IN3 => n354, IN4 => n145, 
                           Q => bdo_out(8));
   U239 : AO222X1 port map( IN1 => n160, IN2 => n364, IN3 => bdi_data(8), IN4 
                           => n155, IN5 => n333, IN6 => n158, Q => n159);
   U247 : AO22X1 port map( IN1 => n166, IN2 => n357, IN3 => n354, IN4 => n149, 
                           Q => bdo_out(6));
   U252 : AO22X1 port map( IN1 => n169, IN2 => n359, IN3 => n354, IN4 => n150, 
                           Q => bdo_out(5));
   U255 : AO221X1 port map( IN1 => ramoutd1(5), IN2 => n302, IN3 => 
                           ramoutd1(37), IN4 => n310, IN5 => n171, Q => n169);
   U257 : AO22X1 port map( IN1 => n205, IN2 => n358, IN3 => n354, IN4 => n152, 
                           Q => bdo_out(4));
   U260 : AO221X1 port map( IN1 => ramoutd1(4), IN2 => n302, IN3 => 
                           ramoutd1(36), IN4 => n310, IN5 => n174, Q => n172);
   U261 : AO22X1 port map( IN1 => ramoutd1(100), IN2 => n314, IN3 => 
                           ramoutd1(68), IN4 => n306, Q => n174);
   U268 : XOR2X1 port map( IN1 => n258, IN2 => n178, Q => n64);
   U269 : AO222X1 port map( IN1 => n333, IN2 => n68, IN3 => cu_cd(7), IN4 => 
                           n179, IN5 => n180, IN6 => bdi_data(31), Q => n178);
   U273 : XOR2X1 port map( IN1 => n163, IN2 => n182, Q => n69);
   U277 : AO22X1 port map( IN1 => n9, IN2 => n359, IN3 => n354, IN4 => n62, Q 
                           => bdo_out(2));
   U283 : XOR2X1 port map( IN1 => n74, IN2 => n187, Q => n72);
   U288 : XOR2X1 port map( IN1 => n7, IN2 => n189, Q => n75);
   U292 : AO22X1 port map( IN1 => n269, IN2 => n357, IN3 => n355, IN4 => n78, Q
                           => bdo_out(27));
   U293 : XOR2X1 port map( IN1 => n269, IN2 => n191, Q => n78);
   U294 : AO222X1 port map( IN1 => n333, IN2 => n80, IN3 => cu_cd(3), IN4 => 
                           n179, IN5 => bdi_data(27), IN6 => n180, Q => n191);
   U297 : AO22X1 port map( IN1 => n273, IN2 => n358, IN3 => n355, IN4 => n81, Q
                           => bdo_out(26));
   U298 : XOR2X1 port map( IN1 => n273, IN2 => n193, Q => n81);
   U303 : XOR2X1 port map( IN1 => n11, IN2 => n195, Q => n84);
   U307 : AO22X1 port map( IN1 => n251, IN2 => n359, IN3 => n355, IN4 => n90, Q
                           => bdo_out(24));
   U308 : XNOR2X1 port map( IN1 => n197, IN2 => n367, Q => n90);
   U309 : AO221X1 port map( IN1 => n333, IN2 => n91, IN3 => bdi_data(24), IN4 
                           => n180, IN5 => n198, Q => n197);
   U311 : AO221X1 port map( IN1 => n302, IN2 => ramoutd1(24), IN3 => 
                           ramoutd1(56), IN4 => n310, IN5 => n199, Q => n91);
   U313 : AO22X1 port map( IN1 => n97, IN2 => n359, IN3 => n355, IN4 => n93, Q 
                           => bdo_out(23));
   U318 : AO22X1 port map( IN1 => n100, IN2 => n357, IN3 => n355, IN4 => n98, Q
                           => bdo_out(22));
   U323 : AO22X1 port map( IN1 => n103, IN2 => n357, IN3 => n355, IN4 => n101, 
                           Q => bdo_out(21));
   U328 : AO22X1 port map( IN1 => n12, IN2 => n357, IN3 => n355, IN4 => n104, Q
                           => bdo_out(20));
   U333 : AO22X1 port map( IN1 => n8, IN2 => n357, IN3 => n355, IN4 => n63, Q 
                           => bdo_out(1));
   U336 : AO221X1 port map( IN1 => n302, IN2 => ramoutd1(1), IN3 => 
                           ramoutd1(33), IN4 => n310, IN5 => n211, Q => n209);
   U338 : AO22X1 port map( IN1 => n109, IN2 => n357, IN3 => n355, IN4 => n107, 
                           Q => bdo_out(19));
   U348 : AO22X1 port map( IN1 => n236, IN2 => n358, IN3 => n355, IN4 => n113, 
                           Q => bdo_out(17));
   U353 : AO22X1 port map( IN1 => n255, IN2 => n358, IN3 => n356, IN4 => n120, 
                           Q => bdo_out(16));
   U354 : XNOR2X1 port map( IN1 => n218, IN2 => n366, Q => n120);
   U355 : AO222X1 port map( IN1 => n117, IN2 => n160, IN3 => bdi_data(16), IN4 
                           => n201, IN5 => n156, IN6 => n121, Q => n218);
   U358 : AO22X1 port map( IN1 => n125, IN2 => n358, IN3 => n356, IN4 => n122, 
                           Q => bdo_out(15));
   U373 : AO22X1 port map( IN1 => n238, IN2 => n359, IN3 => n356, IN4 => n133, 
                           Q => bdo_out(12));
   U378 : AO22X1 port map( IN1 => n220, IN2 => n359, IN3 => n356, IN4 => n136, 
                           Q => bdo_out(11));
   U383 : AO22X1 port map( IN1 => n141, IN2 => n359, IN3 => n356, IN4 => n139, 
                           Q => bdo_out(10));
   U388 : AO22X1 port map( IN1 => n10, IN2 => n359, IN3 => n356, IN4 => n153, Q
                           => bdo_out(0));
   U389 : XOR2X1 port map( IN1 => n233, IN2 => n10, Q => n153);
   U390 : AO222X1 port map( IN1 => n88, IN2 => n160, IN3 => bdi_data(0), IN4 =>
                           n164, IN5 => n156, IN6 => n232, Q => n233);
   U391 : AO21X1 port map( IN1 => n160, IN2 => n364, IN3 => n155, Q => n164);
   U392 : AO21X1 port map( IN1 => n117, IN2 => n160, IN3 => n201, Q => n155);
   U393 : AO21X1 port map( IN1 => n87, IN2 => n160, IN3 => n180, Q => n201);
   U3 : DELLN2X2 port map( INP => ramoutd1(110), Z => n250);
   U4 : AO22X2 port map( IN1 => n112, IN2 => n358, IN3 => n110, IN4 => n355, Q 
                           => bdo_out(18));
   U5 : DELLN2X2 port map( INP => ramoutd1(125), Z => n1);
   U6 : INVX0 port map( INP => n121, ZN => n2);
   U7 : DELLN2X2 port map( INP => ramoutd1(114), Z => n3);
   U8 : AO22X2 port map( IN1 => n74, IN2 => n358, IN3 => n354, IN4 => n72, Q =>
                           bdo_out(29));
   U9 : DELLN2X2 port map( INP => ramoutd1(104), Z => n4);
   U10 : AO22X2 port map( IN1 => ramoutd1(125), IN2 => n314, IN3 => 
                           ramoutd1(93), IN4 => n306, Q => n188);
   U11 : AO221X2 port map( IN1 => ramoutd1(14), IN2 => n302, IN3 => 
                           ramoutd1(46), IN4 => n310, IN5 => n223, Q => n260);
   U12 : AO221X1 port map( IN1 => key(18), IN2 => n337, IN3 => n110, IN4 => 
                           n335, IN5 => n111, Q => n5);
   U13 : DELLN2X2 port map( INP => ramoutd1(122), Z => n6);
   U14 : AO22X2 port map( IN1 => bdi_data(18), IN2 => n95, IN3 => n96, IN4 => 
                           n112, Q => n111);
   U15 : NBUFFX2 port map( INP => n77, Z => n7);
   U16 : NBUFFX2 port map( INP => n209, Z => n8);
   U17 : NBUFFX2 port map( INP => n184, Z => n9);
   U18 : AO22X2 port map( IN1 => ramoutd1(101), IN2 => n314, IN3 => 
                           ramoutd1(69), IN4 => n306, Q => n171);
   U19 : NBUFFX2 port map( INP => n232, Z => n10);
   U20 : AO221X2 port map( IN1 => ramoutd1(22), IN2 => n302, IN3 => 
                           ramoutd1(54), IN4 => n310, IN5 => n204, Q => n100);
   U21 : AO22X2 port map( IN1 => ramoutd1(111), IN2 => n314, IN3 => 
                           ramoutd1(79), IN4 => n306, Q => n221);
   U22 : NBUFFX2 port map( INP => ramoutd1(79), Z => n222);
   U23 : DELLN1X2 port map( INP => ramoutd1(67), Z => n210);
   U24 : AO22X2 port map( IN1 => ramoutd1(99), IN2 => n314, IN3 => ramoutd1(67)
                           , IN4 => n306, Q => n177);
   U25 : NBUFFX2 port map( INP => n86, Z => n11);
   U26 : AO221X1 port map( IN1 => ramoutd1(25), IN2 => n369, IN3 => 
                           ramoutd1(57), IN4 => n310, IN5 => n196, Q => n86);
   U27 : AO22X1 port map( IN1 => n307, IN2 => n35, IN3 => ramoutd1(88), IN4 => 
                           n344, Q => cyc_state_update(88));
   U28 : AO22X2 port map( IN1 => ramoutd1(120), IN2 => n314, IN3 => 
                           ramoutd1(88), IN4 => n306, Q => n199);
   U29 : AO22X2 port map( IN1 => ramoutd1(106), IN2 => n314, IN3 => 
                           ramoutd1(74), IN4 => n306, Q => n231);
   U30 : AO22X2 port map( IN1 => bdi_data(21), IN2 => n95, IN3 => n96, IN4 => 
                           n103, Q => n102);
   U31 : XOR2X1 port map( IN1 => n159, IN2 => n158, Q => n145);
   U32 : AO22X1 port map( IN1 => bdi_data(29), IN2 => n66, IN3 => n67, IN4 => 
                           n74, Q => n73);
   U33 : AO221X2 port map( IN1 => ramoutd1(29), IN2 => n302, IN3 => 
                           ramoutd1(61), IN4 => n310, IN5 => n188, Q => n74);
   U34 : NBUFFX2 port map( INP => n106, Z => n12);
   U35 : NBUFFX2 port map( INP => n144, Z => n13);
   U36 : DELLN2X2 port map( INP => ramoutd1(83), Z => n14);
   U37 : AO22X2 port map( IN1 => ramoutd1(115), IN2 => n350, IN3 => 
                           ramoutd1(83), IN4 => n306, Q => n213);
   U38 : AO22X2 port map( IN1 => bdi_data(28), IN2 => n66, IN3 => n67, IN4 => 
                           n7, Q => n76);
   U39 : AO221X1 port map( IN1 => key(25), IN2 => n338, IN3 => n84, IN4 => n336
                           , IN5 => n85, Q => n15);
   U40 : NAND2X4 port map( IN1 => n37, IN2 => n34, QN => n16);
   U41 : NAND2X0 port map( IN1 => n20, IN2 => n17, QN => n195);
   U42 : INVX4 port map( INP => n16, ZN => n17);
   U43 : NAND2X0 port map( IN1 => bdi_data(25), IN2 => n180, QN => n37);
   U44 : NAND2X0 port map( IN1 => n333, IN2 => n86, QN => n20);
   U45 : NAND2X1 port map( IN1 => cu_cd(1), IN2 => n179, QN => n34);
   U47 : NBUFFX32 port map( INP => n156, Z => n333);
   U48 : AO22X1 port map( IN1 => n311, IN2 => n35, IN3 => ramoutd1(56), IN4 => 
                           n340, Q => cyc_state_update(56));
   U49 : DELLN2X2 port map( INP => ramoutd1(78), Z => n55);
   U50 : MUX41X2 port map( IN1 => ramoutd1(112), IN3 => ramoutd1(80), IN2 => 
                           ramoutd1(48), IN4 => ramoutd1(16), S0 => 
                           dcount_in(0), S1 => dcount_in(1), Q => n121);
   U53 : AO221X1 port map( IN1 => key(30), IN2 => n338, IN3 => n69, IN4 => n336
                           , IN5 => n70, Q => n154);
   U55 : NBUFFX2 port map( INP => n71, Z => n163);
   U56 : AO22X1 port map( IN1 => ramoutd1(98), IN2 => n314, IN3 => ramoutd1(66)
                           , IN4 => n306, Q => n186);
   U57 : NAND2X0 port map( IN1 => n333, IN2 => n77, QN => n167);
   U58 : NAND2X1 port map( IN1 => cu_cd(4), IN2 => n179, QN => n170);
   U59 : NAND2X2 port map( IN1 => bdi_data(28), IN2 => n180, QN => n173);
   U60 : NAND3X0 port map( IN1 => n167, IN2 => n170, IN3 => n173, QN => n189);
   U63 : NOR2X1 port map( IN1 => n372, IN2 => xor_sel(0), QN => n179);
   U64 : NOR2X4 port map( IN1 => xor_sel(0), IN2 => xor_sel(1), QN => n180);
   U65 : DELLN1X2 port map( INP => ramoutd1(91), Z => n270);
   U68 : AO22X1 port map( IN1 => ramoutd1(123), IN2 => n314, IN3 => 
                           ramoutd1(91), IN4 => n306, Q => n192);
   U70 : AO22X2 port map( IN1 => n260, IN2 => n358, IN3 => n356, IN4 => n127, Q
                           => bdo_out(14));
   U71 : AO22X1 port map( IN1 => ramoutd1(121), IN2 => n314, IN3 => 
                           ramoutd1(89), IN4 => n306, Q => n196);
   U72 : AO221X2 port map( IN1 => ramoutd1(21), IN2 => n302, IN3 => 
                           ramoutd1(53), IN4 => n310, IN5 => n206, Q => n103);
   U74 : AO221X1 port map( IN1 => key(28), IN2 => n338, IN3 => n75, IN4 => n336
                           , IN5 => n76, Q => n176);
   U75 : AO22X2 port map( IN1 => ramoutd1(118), IN2 => n314, IN3 => 
                           ramoutd1(86), IN4 => n306, Q => n204);
   U77 : AO22X2 port map( IN1 => n7, IN2 => n359, IN3 => n75, IN4 => n354, Q =>
                           bdo_out(28));
   U78 : AO22X2 port map( IN1 => bdi_data(19), IN2 => n95, IN3 => n96, IN4 => 
                           n109, Q => n108);
   U79 : NBUFFX2 port map( INP => n132, Z => n185);
   U80 : AO221X1 port map( IN1 => ramoutd1(13), IN2 => n302, IN3 => 
                           ramoutd1(45), IN4 => n310, IN5 => n225, Q => n132);
   U81 : AO221X2 port map( IN1 => ramoutd1(19), IN2 => n302, IN3 => 
                           ramoutd1(51), IN4 => n310, IN5 => n213, Q => n109);
   U82 : AO22X2 port map( IN1 => n185, IN2 => n359, IN3 => n356, IN4 => n130, Q
                           => bdo_out(13));
   U83 : AO221X1 port map( IN1 => ramoutd1(10), IN2 => n302, IN3 => 
                           ramoutd1(42), IN4 => n310, IN5 => n231, Q => n141);
   U84 : AO221X1 port map( IN1 => key(10), IN2 => n337, IN3 => n335, IN4 => 
                           n139, IN5 => n140, Q => n190);
   U85 : NAND2X1 port map( IN1 => bdi_data(26), IN2 => n180, QN => n267);
   U86 : AO22X2 port map( IN1 => n11, IN2 => n358, IN3 => n84, IN4 => n355, Q 
                           => bdo_out(25));
   U87 : AO221X1 port map( IN1 => ramoutd1(14), IN2 => n302, IN3 => 
                           ramoutd1(46), IN4 => n310, IN5 => n223, Q => n129);
   U88 : AO221X1 port map( IN1 => ramoutd1(15), IN2 => n302, IN3 => 
                           ramoutd1(47), IN4 => n310, IN5 => n221, Q => n125);
   U89 : AO221X1 port map( IN1 => ramoutd1(0), IN2 => n302, IN3 => ramoutd1(32)
                           , IN4 => n310, IN5 => n234, Q => n232);
   U90 : AO22X1 port map( IN1 => ramoutd1(102), IN2 => n314, IN3 => 
                           ramoutd1(70), IN4 => n306, Q => n168);
   U91 : NOR2X0 port map( IN1 => n372, IN2 => n373, QN => n160);
   U93 : AO221X1 port map( IN1 => ramoutd1(18), IN2 => n302, IN3 => 
                           ramoutd1(50), IN4 => n310, IN5 => n215, Q => n112);
   U94 : AO221X1 port map( IN1 => ramoutd1(20), IN2 => n302, IN3 => 
                           ramoutd1(52), IN4 => n310, IN5 => n208, Q => n106);
   U95 : AO22X1 port map( IN1 => n302, IN2 => n25, IN3 => ramoutd1(0), IN4 => 
                           n353, Q => cyc_state_update(0));
   U96 : AO22X1 port map( IN1 => n304, IN2 => n47, IN3 => ramoutd1(13), IN4 => 
                           n353, Q => cyc_state_update(13));
   U97 : AO22X1 port map( IN1 => n311, IN2 => n25, IN3 => ramoutd1(32), IN4 => 
                           n342, Q => cyc_state_update(32));
   U98 : AO22X1 port map( IN1 => n313, IN2 => n51, IN3 => ramoutd1(38), IN4 => 
                           n342, Q => cyc_state_update(38));
   U99 : AO22X1 port map( IN1 => n312, IN2 => n47, IN3 => ramoutd1(45), IN4 => 
                           n341, Q => cyc_state_update(45));
   U101 : AO22X1 port map( IN1 => n307, IN2 => n24, IN3 => ramoutd1(65), IN4 =>
                           n346, Q => cyc_state_update(65));
   U102 : AO22X1 port map( IN1 => n316, IN2 => n47, IN3 => ramoutd1(109), IN4 
                           => n348, Q => cyc_state_update(109));
   U103 : AND2X1 port map( IN1 => n275, IN2 => n276, Q => n200);
   U105 : AO22X1 port map( IN1 => n313, IN2 => n52, IN3 => ramoutd1(37), IN4 =>
                           n342, Q => cyc_state_update(37));
   U106 : AO22X1 port map( IN1 => n312, IN2 => n39, IN3 => ramoutd1(52), IN4 =>
                           n340, Q => cyc_state_update(52));
   U107 : DELLN2X2 port map( INP => ramoutd1(69), Z => n203);
   U108 : AO22X1 port map( IN1 => ramoutd1(103), IN2 => n314, IN3 => 
                           ramoutd1(71), IN4 => n306, Q => n165);
   U109 : NBUFFX2 port map( INP => n172, Z => n205);
   U110 : DELLN1X2 port map( INP => ramoutd1(68), Z => n207);
   U111 : AO22X2 port map( IN1 => n314, IN2 => n52, IN3 => ramoutd1(101), IN4 
                           => n349, Q => cyc_state_update(101));
   U113 : NBUFFX2 port map( INP => n175, Z => n212);
   U114 : AO22X1 port map( IN1 => n303, IN2 => n23, IN3 => ramoutd1(2), IN4 => 
                           n351, Q => cyc_state_update(2));
   U115 : DELLN2X2 port map( INP => ramoutd1(127), Z => n214);
   U116 : AO221X1 port map( IN1 => key(17), IN2 => n337, IN3 => n335, IN4 => 
                           n113, IN5 => n114, Q => n216);
   U118 : XOR2X1 port map( IN1 => n282, IN2 => n212, Q => n59);
   U120 : AO22X2 port map( IN1 => n212, IN2 => n358, IN3 => n354, IN4 => n59, Q
                           => bdo_out(3));
   U121 : AO22X1 port map( IN1 => n307, IN2 => n53, IN3 => n207, IN4 => n346, Q
                           => cyc_state_update(68));
   U122 : AO22X1 port map( IN1 => ramoutd1(127), IN2 => n314, IN3 => 
                           ramoutd1(95), IN4 => n306, Q => n181);
   U123 : AO221X1 port map( IN1 => key(12), IN2 => n337, IN3 => n133, IN4 => 
                           n335, IN5 => n134, Q => n219);
   U125 : AO22X1 port map( IN1 => n313, IN2 => n53, IN3 => ramoutd1(36), IN4 =>
                           n342, Q => cyc_state_update(36));
   U126 : AO22X1 port map( IN1 => n307, IN2 => n52, IN3 => n203, IN4 => n346, Q
                           => cyc_state_update(69));
   U127 : AO22X1 port map( IN1 => n303, IN2 => n52, IN3 => ramoutd1(5), IN4 => 
                           n351, Q => cyc_state_update(5));
   U128 : NBUFFX2 port map( INP => n138, Z => n220);
   U129 : AO22X1 port map( IN1 => n309, IN2 => n36, IN3 => ramoutd1(87), IN4 =>
                           n344, Q => cyc_state_update(87));
   U130 : AO221X1 port map( IN1 => ramoutd1(11), IN2 => n302, IN3 => 
                           ramoutd1(43), IN4 => n310, IN5 => n229, Q => n138);
   U131 : AO221X1 port map( IN1 => key(15), IN2 => n337, IN3 => n335, IN4 => 
                           n122, IN5 => n123, Q => n224);
   U132 : DELLN2X2 port map( INP => ramoutd1(86), Z => n226);
   U133 : AO221X1 port map( IN1 => key(22), IN2 => n338, IN3 => n98, IN4 => 
                           n335, IN5 => n99, Q => n228);
   U134 : AO221X1 port map( IN1 => key(22), IN2 => n338, IN3 => n98, IN4 => 
                           n335, IN5 => n99, Q => n230);
   U135 : AO221X1 port map( IN1 => key(11), IN2 => n337, IN3 => n136, IN4 => 
                           n335, IN5 => n137, Q => n235);
   U137 : AO22X1 port map( IN1 => n312, IN2 => n235, IN3 => ramoutd1(43), IN4 
                           => n341, Q => cyc_state_update(43));
   U138 : NBUFFX2 port map( INP => n115, Z => n236);
   U139 : DELLN2X2 port map( INP => ramoutd1(119), Z => n237);
   U140 : NBUFFX2 port map( INP => n135, Z => n238);
   U141 : AO221X1 port map( IN1 => ramoutd1(12), IN2 => n302, IN3 => 
                           ramoutd1(44), IN4 => n310, IN5 => n227, Q => n135);
   U142 : AO22X1 port map( IN1 => n315, IN2 => n25, IN3 => ramoutd1(96), IN4 =>
                           n347, Q => cyc_state_update(96));
   U143 : AO221X1 port map( IN1 => ramoutd1(27), IN2 => n302, IN3 => 
                           ramoutd1(59), IN4 => n310, IN5 => n192, Q => n80);
   U144 : AO22X1 port map( IN1 => n303, IN2 => n36, IN3 => ramoutd1(23), IN4 =>
                           n352, Q => cyc_state_update(23));
   U145 : AO22X1 port map( IN1 => n311, IN2 => n36, IN3 => ramoutd1(55), IN4 =>
                           n340, Q => cyc_state_update(55));
   U147 : AO221X1 port map( IN1 => ramoutd1(26), IN2 => n302, IN3 => 
                           ramoutd1(58), IN4 => n310, IN5 => n194, Q => n83);
   U148 : AO221X1 port map( IN1 => key(21), IN2 => n337, IN3 => n101, IN4 => 
                           n335, IN5 => n102, Q => n239);
   U150 : AO221X1 port map( IN1 => key(27), IN2 => n338, IN3 => n78, IN4 => 
                           n336, IN5 => n79, Q => n240);
   U151 : AO22X1 port map( IN1 => n302, IN2 => n51, IN3 => ramoutd1(6), IN4 => 
                           n351, Q => cyc_state_update(6));
   U153 : AO221X1 port map( IN1 => ramoutd1(6), IN2 => n302, IN3 => 
                           ramoutd1(38), IN4 => n310, IN5 => n168, Q => n166);
   U154 : AO22X1 port map( IN1 => n308, IN2 => n224, IN3 => n222, IN4 => n345, 
                           Q => cyc_state_update(79));
   U156 : AO22X1 port map( IN1 => n312, IN2 => n224, IN3 => ramoutd1(47), IN4 
                           => n341, Q => cyc_state_update(47));
   U157 : AO22X1 port map( IN1 => n316, IN2 => n36, IN3 => n237, IN4 => n348, Q
                           => cyc_state_update(119));
   U158 : AO221X1 port map( IN1 => ramoutd1(2), IN2 => n302, IN3 => 
                           ramoutd1(34), IN4 => n310, IN5 => n186, Q => n184);
   U160 : AO22X1 port map( IN1 => n317, IN2 => n49, IN3 => ramoutd1(107), IN4 
                           => n349, Q => cyc_state_update(107));
   U162 : AO22X1 port map( IN1 => n305, IN2 => n235, IN3 => ramoutd1(11), IN4 
                           => n353, Q => cyc_state_update(11));
   U163 : AO221X1 port map( IN1 => key(14), IN2 => n337, IN3 => n335, IN4 => 
                           n127, IN5 => n128, Q => n241);
   U164 : AO22X1 port map( IN1 => n228, IN2 => n311, IN3 => ramoutd1(54), IN4 
                           => n340, Q => cyc_state_update(54));
   U165 : AO22X1 port map( IN1 => n316, IN2 => n228, IN3 => ramoutd1(118), IN4 
                           => n348, Q => cyc_state_update(118));
   U168 : AO22X1 port map( IN1 => n230, IN2 => n309, IN3 => n226, IN4 => n344, 
                           Q => cyc_state_update(86));
   U171 : AO22X1 port map( IN1 => n304, IN2 => n230, IN3 => ramoutd1(22), IN4 
                           => n352, Q => cyc_state_update(22));
   U172 : DELLN2X2 port map( INP => ramoutd1(111), Z => n242);
   U175 : DELLN2X2 port map( INP => ramoutd1(75), Z => n243);
   U176 : AO22X1 port map( IN1 => n312, IN2 => n40, IN3 => ramoutd1(51), IN4 =>
                           n341, Q => cyc_state_update(51));
   U177 : AO221X1 port map( IN1 => ramoutd1(8), IN2 => n302, IN3 => 
                           ramoutd1(40), IN4 => n311, IN5 => n161, Q => n158);
   U180 : AO22X1 port map( IN1 => n42, IN2 => n316, IN3 => ramoutd1(113), IN4 
                           => n348, Q => cyc_state_update(113));
   U183 : DELLN1X2 port map( INP => ramoutd1(100), Z => n321);
   U186 : AO22X1 port map( IN1 => n312, IN2 => n48, IN3 => ramoutd1(44), IN4 =>
                           n341, Q => cyc_state_update(44));
   U187 : AO22X1 port map( IN1 => n304, IN2 => n48, IN3 => ramoutd1(12), IN4 =>
                           n353, Q => cyc_state_update(12));
   U189 : AO221X1 port map( IN1 => key(27), IN2 => n338, IN3 => n78, IN4 => 
                           n336, IN5 => n79, Q => n31);
   U190 : AO22X1 port map( IN1 => n49, IN2 => n308, IN3 => n243, IN4 => n345, Q
                           => cyc_state_update(75));
   U192 : AO22X1 port map( IN1 => n312, IN2 => n5, IN3 => ramoutd1(50), IN4 => 
                           n341, Q => cyc_state_update(50));
   U196 : DELLN2X2 port map( INP => ramoutd1(81), Z => n244);
   U200 : AO22X1 port map( IN1 => n304, IN2 => n39, IN3 => ramoutd1(20), IN4 =>
                           n352, Q => cyc_state_update(20));
   U202 : DELLN2X2 port map( INP => ramoutd1(76), Z => n245);
   U203 : AO22X1 port map( IN1 => n312, IN2 => n21, IN3 => ramoutd1(35), IN4 =>
                           n342, Q => cyc_state_update(35));
   U206 : AO22X1 port map( IN1 => n316, IN2 => n45, IN3 => n242, IN4 => n348, Q
                           => cyc_state_update(111));
   U209 : AO22X1 port map( IN1 => n305, IN2 => n21, IN3 => ramoutd1(3), IN4 => 
                           n351, Q => cyc_state_update(3));
   U212 : AO221X1 port map( IN1 => n334, IN2 => n145, IN3 => 
                           cyc_state_update_sel(1), IN4 => n361, IN5 => n146, Q
                           => n246);
   U215 : AO221X1 port map( IN1 => key(29), IN2 => n338, IN3 => n72, IN4 => 
                           n336, IN5 => n73, Q => n247);
   U224 : AO22X1 port map( IN1 => n32, IN2 => n308, IN3 => ramoutd1(90), IN4 =>
                           n344, Q => cyc_state_update(90));
   U226 : AO22X1 port map( IN1 => n32, IN2 => n316, IN3 => n6, IN4 => n347, Q 
                           => cyc_state_update(122));
   U228 : AO22X1 port map( IN1 => n312, IN2 => n42, IN3 => ramoutd1(49), IN4 =>
                           n341, Q => cyc_state_update(49));
   U230 : AO22X1 port map( IN1 => n307, IN2 => n21, IN3 => n210, IN4 => n346, Q
                           => cyc_state_update(67));
   U233 : AO22X1 port map( IN1 => n306, IN2 => n25, IN3 => ramoutd1(64), IN4 =>
                           n346, Q => cyc_state_update(64));
   U234 : AO22X2 port map( IN1 => ramoutd1(96), IN2 => n314, IN3 => 
                           ramoutd1(64), IN4 => n306, Q => n234);
   U235 : AO22X1 port map( IN1 => n304, IN2 => n24, IN3 => ramoutd1(1), IN4 => 
                           n352, Q => cyc_state_update(1));
   U236 : AO22X1 port map( IN1 => n304, IN2 => n45, IN3 => ramoutd1(15), IN4 =>
                           n353, Q => cyc_state_update(15));
   U238 : AO22X1 port map( IN1 => n308, IN2 => n216, IN3 => n244, IN4 => n345, 
                           Q => cyc_state_update(81));
   U240 : AO22X2 port map( IN1 => ramoutd1(113), IN2 => n314, IN3 => 
                           ramoutd1(81), IN4 => n306, Q => n217);
   U241 : AO22X1 port map( IN1 => n304, IN2 => n216, IN3 => ramoutd1(17), IN4 
                           => n352, Q => cyc_state_update(17));
   U242 : AO221X1 port map( IN1 => ramoutd1(17), IN2 => n302, IN3 => 
                           ramoutd1(49), IN4 => n310, IN5 => n217, Q => n115);
   U243 : AO221X1 port map( IN1 => ramoutd1(30), IN2 => n302, IN3 => 
                           ramoutd1(62), IN4 => n310, IN5 => n183, Q => n71);
   U244 : AO22X1 port map( IN1 => n219, IN2 => n308, IN3 => n245, IN4 => n345, 
                           Q => cyc_state_update(76));
   U245 : AO22X1 port map( IN1 => n307, IN2 => n23, IN3 => ramoutd1(66), IN4 =>
                           n346, Q => cyc_state_update(66));
   U246 : AO22X1 port map( IN1 => n313, IN2 => n23, IN3 => ramoutd1(34), IN4 =>
                           n342, Q => cyc_state_update(34));
   U248 : AO22X1 port map( IN1 => n315, IN2 => n51, IN3 => ramoutd1(102), IN4 
                           => n349, Q => cyc_state_update(102));
   U249 : AO22X1 port map( IN1 => n315, IN2 => n30, IN3 => ramoutd1(124), IN4 
                           => n347, Q => cyc_state_update(124));
   U250 : AO22X1 port map( IN1 => n311, IN2 => n176, IN3 => ramoutd1(60), IN4 
                           => n340, Q => cyc_state_update(60));
   U251 : AO22X1 port map( IN1 => n307, IN2 => n176, IN3 => ramoutd1(92), IN4 
                           => n344, Q => cyc_state_update(92));
   U253 : AO22X1 port map( IN1 => n308, IN2 => n18, IN3 => ramoutd1(73), IN4 =>
                           n345, Q => cyc_state_update(73));
   U254 : AO22X1 port map( IN1 => n316, IN2 => n219, IN3 => ramoutd1(108), IN4 
                           => n348, Q => cyc_state_update(108));
   U256 : AO22X1 port map( IN1 => ramoutd1(108), IN2 => n314, IN3 => 
                           ramoutd1(76), IN4 => n306, Q => n227);
   U258 : DELLN2X2 port map( INP => ramoutd1(9), Z => n248);
   U259 : AO22X1 port map( IN1 => n302, IN2 => n18, IN3 => n248, IN4 => n351, Q
                           => cyc_state_update(9));
   U262 : AO22X1 port map( IN1 => n38, IN2 => n304, IN3 => ramoutd1(21), IN4 =>
                           n352, Q => cyc_state_update(21));
   U263 : AO22X1 port map( IN1 => n308, IN2 => n40, IN3 => n14, IN4 => n345, Q 
                           => cyc_state_update(83));
   U264 : DELLN2X2 port map( INP => ramoutd1(28), Z => n249);
   U265 : AO22X2 port map( IN1 => bdi_data(30), IN2 => n66, IN3 => n67, IN4 => 
                           n163, Q => n70);
   U266 : AO22X2 port map( IN1 => n163, IN2 => n359, IN3 => n69, IN4 => n354, Q
                           => bdo_out(30));
   U267 : AO22X1 port map( IN1 => n30, IN2 => n303, IN3 => n249, IN4 => n351, Q
                           => cyc_state_update(28));
   U270 : AO22X1 port map( IN1 => n315, IN2 => n31, IN3 => ramoutd1(123), IN4 
                           => n347, Q => cyc_state_update(123));
   U271 : AO22X1 port map( IN1 => n311, IN2 => n240, IN3 => ramoutd1(59), IN4 
                           => n340, Q => cyc_state_update(59));
   U272 : AO22X1 port map( IN1 => n316, IN2 => n41, IN3 => n3, IN4 => n348, Q 
                           => cyc_state_update(114));
   U274 : AO22X1 port map( IN1 => n303, IN2 => n240, IN3 => ramoutd1(27), IN4 
                           => n352, Q => cyc_state_update(27));
   U275 : AO22X1 port map( IN1 => n304, IN2 => n5, IN3 => ramoutd1(18), IN4 => 
                           n352, Q => cyc_state_update(18));
   U276 : AO22X1 port map( IN1 => n311, IN2 => n32, IN3 => ramoutd1(58), IN4 =>
                           n340, Q => cyc_state_update(58));
   U278 : AO22X1 port map( IN1 => n303, IN2 => n32, IN3 => ramoutd1(26), IN4 =>
                           n352, Q => cyc_state_update(26));
   U279 : AO22X1 port map( IN1 => n307, IN2 => n51, IN3 => ramoutd1(70), IN4 =>
                           n346, Q => cyc_state_update(70));
   U280 : AO22X1 port map( IN1 => n311, IN2 => n38, IN3 => ramoutd1(53), IN4 =>
                           n340, Q => cyc_state_update(53));
   U281 : IBUFFX16 port map( INP => n367, ZN => n251);
   U282 : DELLN2X2 port map( INP => ramoutd1(82), Z => n252);
   U284 : AO22X1 port map( IN1 => n308, IN2 => n41, IN3 => n252, IN4 => n345, Q
                           => cyc_state_update(82));
   U285 : AO22X1 port map( IN1 => n47, IN2 => n308, IN3 => ramoutd1(77), IN4 =>
                           n345, Q => cyc_state_update(77));
   U286 : DELLN1X2 port map( INP => ramoutd1(117), Z => n318);
   U287 : AO222X1 port map( IN1 => key(24), IN2 => n338, IN3 => n360, IN4 => 
                           n89, IN5 => n334, IN6 => n90, Q => n253);
   U289 : DELLN2X2 port map( INP => ramoutd1(95), Z => n254);
   U290 : AO22X2 port map( IN1 => n258, IN2 => n358, IN3 => n64, IN4 => n354, Q
                           => bdo_out(31));
   U291 : AO22X1 port map( IN1 => n29, IN2 => n315, IN3 => n1, IN4 => n347, Q 
                           => cyc_state_update(125));
   U295 : AO22X1 port map( IN1 => n314, IN2 => ramoutd1(104), IN3 => 
                           ramoutd1(72), IN4 => n306, Q => n161);
   U296 : AO22X1 port map( IN1 => n311, IN2 => n247, IN3 => ramoutd1(61), IN4 
                           => n340, Q => cyc_state_update(61));
   U299 : AO22X1 port map( IN1 => n29, IN2 => n303, IN3 => ramoutd1(29), IN4 =>
                           n351, Q => cyc_state_update(29));
   U300 : AO22X1 port map( IN1 => n317, IN2 => n18, IN3 => ramoutd1(105), IN4 
                           => n349, Q => cyc_state_update(105));
   U301 : AO221X1 port map( IN1 => ramoutd1(73), IN2 => n306, IN3 => 
                           ramoutd1(105), IN4 => n314, IN5 => n157, Q => n144);
   U302 : AO22X1 port map( IN1 => n315, IN2 => n154, IN3 => ramoutd1(126), IN4 
                           => n347, Q => cyc_state_update(126));
   U304 : AO22X1 port map( IN1 => n311, IN2 => n28, IN3 => ramoutd1(62), IN4 =>
                           n340, Q => cyc_state_update(62));
   U305 : AO22X1 port map( IN1 => n303, IN2 => n154, IN3 => ramoutd1(30), IN4 
                           => n351, Q => cyc_state_update(30));
   U306 : AO22X2 port map( IN1 => n327, IN2 => n358, IN3 => n354, IN4 => n148, 
                           Q => bdo_out(7));
   U310 : AO22X1 port map( IN1 => n315, IN2 => n23, IN3 => ramoutd1(98), IN4 =>
                           n347, Q => cyc_state_update(98));
   U312 : MUX41X1 port map( IN1 => ramoutd1(124), IN3 => ramoutd1(92), IN2 => 
                           ramoutd1(60), IN4 => ramoutd1(28), S0 => 
                           dcount_in(0), S1 => dcount_in(1), Q => n77);
   U314 : AO22X1 port map( IN1 => n304, IN2 => n40, IN3 => ramoutd1(19), IN4 =>
                           n352, Q => cyc_state_update(19));
   U315 : AO22X1 port map( IN1 => n303, IN2 => n253, IN3 => ramoutd1(24), IN4 
                           => n352, Q => cyc_state_update(24));
   U316 : AO22X1 port map( IN1 => n315, IN2 => n24, IN3 => n256, IN4 => n347, Q
                           => cyc_state_update(97));
   U317 : AO22X1 port map( IN1 => n312, IN2 => n43, IN3 => ramoutd1(48), IN4 =>
                           n341, Q => cyc_state_update(48));
   U319 : AO22X1 port map( IN1 => n315, IN2 => n253, IN3 => ramoutd1(120), IN4 
                           => n347, Q => cyc_state_update(120));
   U320 : AO22X1 port map( IN1 => n312, IN2 => n50, IN3 => ramoutd1(42), IN4 =>
                           n341, Q => cyc_state_update(42));
   U321 : AO22X1 port map( IN1 => n317, IN2 => n50, IN3 => ramoutd1(106), IN4 
                           => n349, Q => cyc_state_update(106));
   U322 : AO22X1 port map( IN1 => n305, IN2 => n50, IN3 => ramoutd1(10), IN4 =>
                           n353, Q => cyc_state_update(10));
   U324 : INVX0 port map( INP => n2, ZN => n255);
   U325 : DELLN2X2 port map( INP => ramoutd1(97), Z => n256);
   U326 : INVX0 port map( INP => n68, ZN => n257);
   U327 : INVX0 port map( INP => n257, ZN => n258);
   U329 : AO221X1 port map( IN1 => ramoutd1(31), IN2 => n302, IN3 => 
                           ramoutd1(63), IN4 => n310, IN5 => n181, Q => n68);
   U330 : AO22X1 port map( IN1 => n314, IN2 => ramoutd1(97), IN3 => 
                           ramoutd1(65), IN4 => n306, Q => n211);
   U331 : AO221X1 port map( IN1 => key(31), IN2 => n338, IN3 => n64, IN4 => 
                           n334, IN5 => n65, Q => n259);
   U332 : AO221X1 port map( IN1 => key(14), IN2 => n337, IN3 => n335, IN4 => 
                           n127, IN5 => n128, Q => n46);
   U334 : AO22X1 port map( IN1 => n307, IN2 => n33, IN3 => ramoutd1(72), IN4 =>
                           n345, Q => cyc_state_update(72));
   U335 : AO22X1 port map( IN1 => n246, IN2 => n312, IN3 => ramoutd1(40), IN4 
                           => n341, Q => cyc_state_update(40));
   U337 : AO22X1 port map( IN1 => n302, IN2 => n33, IN3 => ramoutd1(8), IN4 => 
                           n351, Q => cyc_state_update(8));
   U339 : AO22X1 port map( IN1 => n303, IN2 => n26, IN3 => ramoutd1(31), IN4 =>
                           n351, Q => cyc_state_update(31));
   U340 : AO22X1 port map( IN1 => n306, IN2 => n26, IN3 => n254, IN4 => n344, Q
                           => cyc_state_update(95));
   U341 : AO22X1 port map( IN1 => n311, IN2 => n259, IN3 => ramoutd1(63), IN4 
                           => n340, Q => cyc_state_update(63));
   U342 : AO22X1 port map( IN1 => n259, IN2 => n315, IN3 => n214, IN4 => n347, 
                           Q => cyc_state_update(127));
   U343 : DELLN2X2 port map( INP => ramoutd1(71), Z => n261);
   U344 : AO22X2 port map( IN1 => ramoutd1(107), IN2 => n314, IN3 => 
                           ramoutd1(75), IN4 => n306, Q => n229);
   U345 : AO22X1 port map( IN1 => n314, IN2 => ramoutd1(126), IN3 => 
                           ramoutd1(94), IN4 => n306, Q => n183);
   U346 : AO221X1 port map( IN1 => n302, IN2 => ramoutd1(23), IN3 => 
                           ramoutd1(55), IN4 => n310, IN5 => n202, Q => n97);
   U347 : AO22X1 port map( IN1 => n304, IN2 => n43, IN3 => ramoutd1(16), IN4 =>
                           n353, Q => cyc_state_update(16));
   U349 : AO22X1 port map( IN1 => ramoutd1(117), IN2 => n314, IN3 => 
                           ramoutd1(85), IN4 => n306, Q => n206);
   U350 : AO22X1 port map( IN1 => n315, IN2 => n15, IN3 => ramoutd1(121), IN4 
                           => n347, Q => cyc_state_update(121));
   U351 : AO22X1 port map( IN1 => n303, IN2 => n15, IN3 => ramoutd1(25), IN4 =>
                           n352, Q => cyc_state_update(25));
   U352 : AO22X1 port map( IN1 => n314, IN2 => ramoutd1(116), IN3 => 
                           ramoutd1(84), IN4 => n306, Q => n208);
   U356 : AO221X1 port map( IN1 => ramoutd1(3), IN2 => n302, IN3 => 
                           ramoutd1(35), IN4 => n310, IN5 => n177, Q => n175);
   U357 : AO22X1 port map( IN1 => n304, IN2 => n46, IN3 => ramoutd1(14), IN4 =>
                           n353, Q => cyc_state_update(14));
   U359 : XOR2X1 port map( IN1 => n283, IN2 => n9, Q => n62);
   U360 : INVX0 port map( INP => n367, ZN => n264);
   U361 : AO22X2 port map( IN1 => ramoutd1(114), IN2 => n314, IN3 => 
                           ramoutd1(82), IN4 => n306, Q => n215);
   U362 : AO22X2 port map( IN1 => n312, IN2 => n18, IN3 => ramoutd1(41), IN4 =>
                           n341, Q => cyc_state_update(41));
   U363 : AO22X1 port map( IN1 => ramoutd1(41), IN2 => n311, IN3 => n302, IN4 
                           => ramoutd1(9), Q => n157);
   U364 : DELLN2X2 port map( INP => ramoutd1(99), Z => n325);
   U365 : AO22X2 port map( IN1 => ramoutd1(122), IN2 => n314, IN3 => 
                           ramoutd1(90), IN4 => n306, Q => n194);
   U366 : AO22X1 port map( IN1 => ramoutd1(119), IN2 => n314, IN3 => 
                           ramoutd1(87), IN4 => n306, Q => n202);
   U367 : AO221X1 port map( IN1 => ramoutd1(7), IN2 => n302, IN3 => 
                           ramoutd1(39), IN4 => n311, IN5 => n165, Q => n162);
   U368 : DELLN2X2 port map( INP => ramoutd1(4), Z => n319);
   U369 : AO22X1 port map( IN1 => n314, IN2 => ramoutd1(110), IN3 => 
                           ramoutd1(78), IN4 => n306, Q => n223);
   U370 : DELLN2X2 port map( INP => ramoutd1(115), Z => n262);
   U371 : IBUFFX16 port map( INP => n368, ZN => n263);
   U372 : NAND2X0 port map( IN1 => n333, IN2 => n83, QN => n265);
   U374 : NAND2X1 port map( IN1 => cu_cd(2), IN2 => n179, QN => n266);
   U375 : NAND3X0 port map( IN1 => n265, IN2 => n266, IN3 => n267, QN => n193);
   U376 : INVX0 port map( INP => n80, ZN => n268);
   U377 : INVX0 port map( INP => n268, ZN => n269);
   U379 : DELLN2X2 port map( INP => ramoutd1(89), Z => n271);
   U380 : XOR2X1 port map( IN1 => n12, IN2 => n291, Q => n104);
   U381 : INVX0 port map( INP => n83, ZN => n272);
   U382 : INVX0 port map( INP => n272, ZN => n273);
   U384 : AO22X2 port map( IN1 => bdi_data(17), IN2 => n95, IN3 => n96, IN4 => 
                           n236, Q => n114);
   U385 : NAND2X0 port map( IN1 => n274, IN2 => n200, QN => n182);
   U386 : NAND2X0 port map( IN1 => n156, IN2 => n71, QN => n274);
   U387 : NAND2X1 port map( IN1 => cu_cd(6), IN2 => n179, QN => n275);
   U394 : NAND2X0 port map( IN1 => bdi_data(30), IN2 => n180, QN => n276);
   U395 : AO22X2 port map( IN1 => bdi_data(31), IN2 => n66, IN3 => n67, IN4 => 
                           n258, Q => n65);
   U396 : NAND2X0 port map( IN1 => n333, IN2 => n74, QN => n277);
   U397 : NAND2X1 port map( IN1 => cu_cd(5), IN2 => n179, QN => n278);
   U398 : NAND2X0 port map( IN1 => bdi_data(29), IN2 => n180, QN => n279);
   U399 : NAND3X0 port map( IN1 => n277, IN2 => n278, IN3 => n279, QN => n187);
   U400 : DELLN2X2 port map( INP => ramoutd1(103), Z => n326);
   U401 : DELLN2X2 port map( INP => ramoutd1(93), Z => n280);
   U402 : XOR2X1 port map( IN1 => n220, IN2 => n288, Q => n136);
   U403 : AO22X2 port map( IN1 => bdi_data(25), IN2 => n66, IN3 => n67, IN4 => 
                           n11, Q => n85);
   U404 : AO22X2 port map( IN1 => bdi_data(20), IN2 => n95, IN3 => n96, IN4 => 
                           n12, Q => n105);
   U405 : AO22X2 port map( IN1 => bdi_data(26), IN2 => n66, IN3 => n67, IN4 => 
                           n273, Q => n82);
   U406 : INVX0 port map( INP => n92, ZN => n363);
   U407 : INVX0 port map( INP => n118, ZN => n362);
   U408 : INVX0 port map( INP => n357, ZN => n354);
   U409 : INVX0 port map( INP => n357, ZN => n355);
   U410 : INVX0 port map( INP => n359, ZN => n356);
   U411 : NBUFFX2 port map( INP => n156, Z => n332);
   U412 : INVX0 port map( INP => xor_sel(0), ZN => n373);
   U413 : INVX0 port map( INP => n116, ZN => n360);
   U414 : NOR2X0 port map( IN1 => n116, IN2 => n92, QN => n96);
   U415 : NOR2X0 port map( IN1 => n116, IN2 => n118, QN => n95);
   U416 : NBUFFX2 port map( INP => n58, Z => n334);
   U417 : NBUFFX2 port map( INP => n58, Z => n335);
   U418 : NBUFFX2 port map( INP => n57, Z => n337);
   U419 : NBUFFX2 port map( INP => n57, Z => n338);
   U420 : NBUFFX2 port map( INP => n58, Z => n336);
   U421 : NBUFFX2 port map( INP => n57, Z => n339);
   U422 : INVX0 port map( INP => xor_sel(1), ZN => n372);
   U423 : INVX0 port map( INP => extract_sel, ZN => n357);
   U424 : INVX0 port map( INP => extract_sel, ZN => n359);
   U425 : INVX0 port map( INP => extract_sel, ZN => n358);
   U426 : NOR2X0 port map( IN1 => n373, IN2 => xor_sel(1), QN => n156);
   U427 : NBUFFX2 port map( INP => n331, Z => n307);
   U428 : NBUFFX2 port map( INP => n329, Z => n304);
   U429 : NBUFFX2 port map( INP => n329, Z => n303);
   U430 : NBUFFX2 port map( INP => n331, Z => n308);
   U431 : NBUFFX2 port map( INP => n331, Z => n309);
   U432 : NBUFFX2 port map( INP => n329, Z => n305);
   U433 : INVX0 port map( INP => n121, ZN => n366);
   U434 : INVX0 port map( INP => n158, ZN => n368);
   U435 : INVX0 port map( INP => n91, ZN => n367);
   U436 : NAND2X0 port map( IN1 => cyc_state_update_sel(1), IN2 => 
                           cyc_state_update_sel(0), QN => n116);
   U437 : NOR2X0 port map( IN1 => n361, IN2 => cyc_state_update_sel(1), QN => 
                           n57);
   U438 : NOR2X0 port map( IN1 => cyc_state_update_sel(0), IN2 => 
                           cyc_state_update_sel(1), QN => n58);
   U439 : INVX0 port map( INP => cyc_state_update_sel(0), ZN => n361);
   U440 : NBUFFX2 port map( INP => n343, Z => n311);
   U441 : NOR2X0 port map( IN1 => n314, IN2 => n306, QN => n60);
   U442 : NOR2X0 port map( IN1 => n310, IN2 => n302, QN => n54);
   U443 : NBUFFX2 port map( INP => n328, Z => n302);
   U444 : NBUFFX2 port map( INP => n369, Z => n328);
   U445 : NBUFFX2 port map( INP => n330, Z => n306);
   U446 : NBUFFX2 port map( INP => n370, Z => n330);
   U447 : NBUFFX2 port map( INP => n22, Z => n348);
   U448 : NBUFFX2 port map( INP => n19, Z => n351);
   U449 : NBUFFX2 port map( INP => n19, Z => n352);
   U450 : NBUFFX2 port map( INP => n27, Z => n345);
   U451 : NBUFFX2 port map( INP => n56, Z => n341);
   U452 : NBUFFX2 port map( INP => n56, Z => n340);
   U453 : NBUFFX2 port map( INP => n27, Z => n344);
   U454 : NBUFFX2 port map( INP => n22, Z => n347);
   U455 : NBUFFX2 port map( INP => n56, Z => n342);
   U456 : NBUFFX2 port map( INP => n19, Z => n353);
   U457 : NBUFFX2 port map( INP => n27, Z => n346);
   U458 : NBUFFX2 port map( INP => n22, Z => n349);
   U459 : NBUFFX2 port map( INP => n310, Z => n312);
   U460 : NBUFFX2 port map( INP => n314, Z => n315);
   U461 : NBUFFX2 port map( INP => n314, Z => n316);
   U462 : NBUFFX2 port map( INP => n343, Z => n313);
   U463 : NBUFFX2 port map( INP => n314, Z => n317);
   U464 : NBUFFX2 port map( INP => n369, Z => n329);
   U465 : NBUFFX2 port map( INP => n370, Z => n331);
   U466 : AO22X1 port map( IN1 => n15, IN2 => n307, IN3 => n271, IN4 => n344, Q
                           => cyc_state_update(89));
   U467 : AO22X1 port map( IN1 => n314, IN2 => n53, IN3 => n321, IN4 => n349, Q
                           => cyc_state_update(100));
   U468 : NBUFFX2 port map( INP => n350, Z => n314);
   U469 : INVX0 port map( INP => n300, ZN => n350);
   U470 : NBUFFX2 port map( INP => n343, Z => n310);
   U471 : INVX0 port map( INP => n301, ZN => n343);
   U472 : NAND2X0 port map( IN1 => n54, IN2 => n151, QN => n22);
   U473 : NAND2X0 port map( IN1 => n60, IN2 => n61, QN => n56);
   U474 : NAND2X1 port map( IN1 => n60, IN2 => n301, QN => n19);
   U475 : NAND2X1 port map( IN1 => n54, IN2 => n300, QN => n27);
   U476 : INVX0 port map( INP => n151, ZN => n370);
   U477 : INVX0 port map( INP => n61, ZN => n369);
   U478 : XOR2X1 port map( IN1 => n281, IN2 => n97, Q => n93);
   U479 : AO22X1 port map( IN1 => n201, IN2 => bdi_data(23), IN3 => n332, IN4 
                           => n97, Q => n281);
   U480 : AO22X1 port map( IN1 => cu_cd(0), IN2 => n179, IN3 => n87, IN4 => 
                           n160, Q => n198);
   U481 : AO22X1 port map( IN1 => n164, IN2 => bdi_data(3), IN3 => n175, IN4 =>
                           n332, Q => n282);
   U482 : AO22X1 port map( IN1 => n164, IN2 => bdi_data(2), IN3 => n184, IN4 =>
                           n332, Q => n283);
   U483 : XOR2X1 port map( IN1 => n205, IN2 => n284, Q => n152);
   U484 : AO22X1 port map( IN1 => n164, IN2 => bdi_data(4), IN3 => n332, IN4 =>
                           n172, Q => n284);
   U485 : XOR2X1 port map( IN1 => n8, IN2 => n285, Q => n63);
   U486 : AO22X1 port map( IN1 => n164, IN2 => bdi_data(1), IN3 => n209, IN4 =>
                           n332, Q => n285);
   U487 : XOR2X1 port map( IN1 => n286, IN2 => n327, Q => n148);
   U488 : AO22X1 port map( IN1 => n164, IN2 => bdi_data(7), IN3 => n333, IN4 =>
                           n162, Q => n286);
   U489 : XOR2X1 port map( IN1 => n236, IN2 => n287, Q => n113);
   U490 : AO22X1 port map( IN1 => n201, IN2 => bdi_data(17), IN3 => n115, IN4 
                           => n332, Q => n287);
   U491 : AO22X1 port map( IN1 => n155, IN2 => bdi_data(11), IN3 => n138, IN4 
                           => n332, Q => n288);
   U492 : XOR2X1 port map( IN1 => n103, IN2 => n289, Q => n101);
   U493 : AO22X1 port map( IN1 => n201, IN2 => bdi_data(21), IN3 => n103, IN4 
                           => n332, Q => n289);
   U494 : XOR2X1 port map( IN1 => n290, IN2 => n109, Q => n107);
   U495 : AO22X1 port map( IN1 => n201, IN2 => bdi_data(19), IN3 => n109, IN4 
                           => n332, Q => n290);
   U496 : AO22X1 port map( IN1 => n201, IN2 => bdi_data(20), IN3 => n106, IN4 
                           => n332, Q => n291);
   U497 : XOR2X1 port map( IN1 => n292, IN2 => n112, Q => n110);
   U498 : AO22X1 port map( IN1 => n201, IN2 => bdi_data(18), IN3 => n332, IN4 
                           => n112, Q => n292);
   U499 : XOR2X1 port map( IN1 => n185, IN2 => n293, Q => n130);
   U500 : AO22X1 port map( IN1 => n155, IN2 => bdi_data(13), IN3 => n333, IN4 
                           => n132, Q => n293);
   U501 : XOR2X1 port map( IN1 => n238, IN2 => n294, Q => n133);
   U502 : AO22X1 port map( IN1 => n155, IN2 => bdi_data(12), IN3 => n332, IN4 
                           => n135, Q => n294);
   U503 : XOR2X1 port map( IN1 => n295, IN2 => n260, Q => n127);
   U504 : AO22X1 port map( IN1 => n155, IN2 => bdi_data(14), IN3 => n332, IN4 
                           => n129, Q => n295);
   U505 : XOR2X1 port map( IN1 => n125, IN2 => n296, Q => n122);
   U506 : AO22X1 port map( IN1 => n155, IN2 => bdi_data(15), IN3 => n125, IN4 
                           => n332, Q => n296);
   U507 : XOR2X1 port map( IN1 => n141, IN2 => n297, Q => n139);
   U508 : AO22X1 port map( IN1 => n155, IN2 => bdi_data(10), IN3 => n141, IN4 
                           => n332, Q => n297);
   U509 : XOR2X1 port map( IN1 => n100, IN2 => n298, Q => n98);
   U510 : AO22X1 port map( IN1 => n201, IN2 => bdi_data(22), IN3 => n100, IN4 
                           => n332, Q => n298);
   U511 : XOR2X1 port map( IN1 => n13, IN2 => n299, Q => n142);
   U512 : AO22X1 port map( IN1 => n155, IN2 => bdi_data(9), IN3 => n156, IN4 =>
                           n144, Q => n299);
   U513 : AO22X1 port map( IN1 => bdi_data(22), IN2 => n95, IN3 => n96, IN4 => 
                           n100, Q => n99);
   U514 : OR2X1 port map( IN1 => dcount_in(0), IN2 => dcount_in(1), Q => n300);
   U515 : OR2X1 port map( IN1 => n371, IN2 => dcount_in(0), Q => n301);
   U516 : NAND2X0 port map( IN1 => dcount_in(0), IN2 => n371, QN => n151);
   U517 : NAND2X0 port map( IN1 => dcount_in(0), IN2 => dcount_in(1), QN => n61
                           );
   U518 : INVX0 port map( INP => dcount_in(1), ZN => n371);
   U519 : NOR2X0 port map( IN1 => n87, IN2 => n88, QN => n118);
   U520 : XOR2X1 port map( IN1 => n166, IN2 => n320, Q => n149);
   U521 : AO22X1 port map( IN1 => n164, IN2 => bdi_data(6), IN3 => n166, IN4 =>
                           n333, Q => n320);
   U522 : NAND2X0 port map( IN1 => n314, IN2 => ramoutd1(109), QN => n322);
   U523 : NAND2X0 port map( IN1 => n306, IN2 => ramoutd1(77), QN => n323);
   U524 : NAND2X0 port map( IN1 => n322, IN2 => n323, QN => n225);
   U525 : XOR2X1 port map( IN1 => n169, IN2 => n324, Q => n150);
   U526 : AO22X1 port map( IN1 => n164, IN2 => bdi_data(5), IN3 => n332, IN4 =>
                           n169, Q => n324);
   U527 : NBUFFX2 port map( INP => n162, Z => n327);
   U528 : AND2X1 port map( IN1 => cycd_sel(0), IN2 => cycd_sel(1), Q => n87);
   U529 : INVX0 port map( INP => cycd_sel(1), ZN => n365);
   U530 : NOR2X0 port map( IN1 => n147, IN2 => n116, QN => n124);
   U531 : NOR2X0 port map( IN1 => n364, IN2 => n117, QN => n92);
   U532 : NOR2X0 port map( IN1 => cycd_sel(0), IN2 => cycd_sel(1), QN => n88);
   U533 : INVX0 port map( INP => n147, ZN => n364);
   U534 : NAND2X0 port map( IN1 => cycd_sel(0), IN2 => n365, QN => n147);
   U535 : NOR2X0 port map( IN1 => n365, IN2 => cycd_sel(0), QN => n117);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_LWC_1.all;

entity counter_num_bits5_1 is

   port( clk, load, enable : in std_logic;  start_value : in std_logic_vector 
         (4 downto 0);  q : out std_logic_vector (4 downto 0));

end counter_num_bits5_1;

architecture SYN_Behavioral of counter_num_bits5_1 is

   component XOR2X1
      port( IN1, IN2 : in std_logic;  Q : out std_logic);
   end component;
   
   component NOR2X0
      port( IN1, IN2 : in std_logic;  QN : out std_logic);
   end component;
   
   component HADDX1
      port( A0, B0 : in std_logic;  C1, SO : out std_logic);
   end component;
   
   component AO222X1
      port( IN1, IN2, IN3, IN4, IN5, IN6 : in std_logic;  Q : out std_logic);
   end component;
   
   component DFFX1
      port( D, CLK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal q_4_port, q_3_port, q_2_port, q_1_port, q_0_port, N5, N6, N7, N8, n1,
      n2, n3, n4, n5_port, n6_port, n7_port, add_40_carry_2_port, 
      add_40_carry_3_port, add_40_carry_4_port, n8_port, n_1023, n_1024, n_1025
      , n_1026 : std_logic;

begin
   q <= ( q_4_port, q_3_port, q_2_port, q_1_port, q_0_port );
   
   count_reg_0_inst : DFFX1 port map( D => n7_port, CLK => clk, Q => q_0_port, 
                           QN => n8_port);
   count_reg_1_inst : DFFX1 port map( D => n6_port, CLK => clk, Q => q_1_port, 
                           QN => n_1023);
   count_reg_2_inst : DFFX1 port map( D => n5_port, CLK => clk, Q => q_2_port, 
                           QN => n_1024);
   count_reg_3_inst : DFFX1 port map( D => n4, CLK => clk, Q => q_3_port, QN =>
                           n_1025);
   count_reg_4_inst : DFFX1 port map( D => n3, CLK => clk, Q => q_4_port, QN =>
                           n_1026);
   U5 : AO222X1 port map( IN1 => start_value(4), IN2 => load, IN3 => N8, IN4 =>
                           n1, IN5 => q_4_port, IN6 => n2, Q => n3);
   U6 : AO222X1 port map( IN1 => start_value(3), IN2 => load, IN3 => N7, IN4 =>
                           n1, IN5 => q_3_port, IN6 => n2, Q => n4);
   U7 : AO222X1 port map( IN1 => start_value(2), IN2 => load, IN3 => N6, IN4 =>
                           n1, IN5 => q_2_port, IN6 => n2, Q => n5_port);
   U8 : AO222X1 port map( IN1 => start_value(1), IN2 => load, IN3 => N5, IN4 =>
                           n1, IN5 => q_1_port, IN6 => n2, Q => n6_port);
   U9 : AO222X1 port map( IN1 => start_value(0), IN2 => load, IN3 => n8_port, 
                           IN4 => n1, IN5 => q_0_port, IN6 => n2, Q => n7_port)
                           ;
   add_40_U1_1_1 : HADDX1 port map( A0 => q_1_port, B0 => q_0_port, C1 => 
                           add_40_carry_2_port, SO => N5);
   add_40_U1_1_2 : HADDX1 port map( A0 => q_2_port, B0 => add_40_carry_2_port, 
                           C1 => add_40_carry_3_port, SO => N6);
   add_40_U1_1_3 : HADDX1 port map( A0 => q_3_port, B0 => add_40_carry_3_port, 
                           C1 => add_40_carry_4_port, SO => N7);
   U3 : NOR2X0 port map( IN1 => enable, IN2 => load, QN => n2);
   U4 : NOR2X0 port map( IN1 => n2, IN2 => load, QN => n1);
   U10 : XOR2X1 port map( IN1 => add_40_carry_4_port, IN2 => q_4_port, Q => N8)
                           ;

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_LWC_1.all;

entity counter_num_bits4_1_0 is

   port( clk, load, enable : in std_logic;  start_value : in std_logic_vector 
         (3 downto 0);  q : out std_logic_vector (3 downto 0));

end counter_num_bits4_1_0;

architecture SYN_Behavioral of counter_num_bits4_1_0 is

   component NOR2X0
      port( IN1, IN2 : in std_logic;  QN : out std_logic);
   end component;
   
   component NOR4X0
      port( IN1, IN2, IN3, IN4 : in std_logic;  QN : out std_logic);
   end component;
   
   component INVX0
      port( INP : in std_logic;  ZN : out std_logic);
   end component;
   
   component AO222X1
      port( IN1, IN2, IN3, IN4, IN5, IN6 : in std_logic;  Q : out std_logic);
   end component;
   
   component NAND3X0
      port( IN1, IN2, IN3 : in std_logic;  QN : out std_logic);
   end component;
   
   component OAI21X1
      port( IN1, IN2, IN3 : in std_logic;  QN : out std_logic);
   end component;
   
   component AO21X1
      port( IN1, IN2, IN3 : in std_logic;  Q : out std_logic);
   end component;
   
   component AO221X1
      port( IN1, IN2, IN3, IN4, IN5 : in std_logic;  Q : out std_logic);
   end component;
   
   component DFFX1
      port( D, CLK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal q_3_port, q_2_port, q_1_port, q_0_port, n1, n2, n6, n7, n8, n9, n10, 
      n11, n12, n13, n14, n15, n16, n17, n3, n4, n5, n_1027, n_1028 : std_logic
      ;

begin
   q <= ( q_3_port, q_2_port, q_1_port, q_0_port );
   
   count_reg_0_inst : DFFX1 port map( D => n17, CLK => clk, Q => q_0_port, QN 
                           => n_1027);
   count_reg_1_inst : DFFX1 port map( D => n16, CLK => clk, Q => q_1_port, QN 
                           => n2);
   count_reg_2_inst : DFFX1 port map( D => n15, CLK => clk, Q => q_2_port, QN 
                           => n1);
   count_reg_3_inst : DFFX1 port map( D => n14, CLK => clk, Q => q_3_port, QN 
                           => n_1028);
   U10 : AO221X1 port map( IN1 => q_3_port, IN2 => n6, IN3 => start_value(3), 
                           IN4 => load, IN5 => n7, Q => n14);
   U11 : AO21X1 port map( IN1 => n5, IN2 => n1, IN3 => n9, Q => n6);
   U12 : AO222X1 port map( IN1 => start_value(2), IN2 => load, IN3 => n10, IN4 
                           => q_1_port, IN5 => q_2_port, IN6 => n9, Q => n15);
   U13 : AO21X1 port map( IN1 => n5, IN2 => n2, IN3 => n11, Q => n9);
   U14 : AO222X1 port map( IN1 => n3, IN2 => n2, IN3 => start_value(1), IN4 => 
                           load, IN5 => q_1_port, IN6 => n11, Q => n16);
   U15 : OAI21X1 port map( IN1 => load, IN2 => q_0_port, IN3 => n4, QN => n11);
   U16 : NAND3X0 port map( IN1 => n4, IN2 => n5, IN3 => q_0_port, QN => n8);
   U17 : AO222X1 port map( IN1 => start_value(0), IN2 => load, IN3 => n12, IN4 
                           => n4, IN5 => n13, IN6 => q_0_port, Q => n17);
   U3 : INVX0 port map( INP => n13, ZN => n4);
   U4 : INVX0 port map( INP => load, ZN => n5);
   U5 : NOR2X0 port map( IN1 => enable, IN2 => load, QN => n13);
   U6 : INVX0 port map( INP => n8, ZN => n3);
   U7 : NOR2X0 port map( IN1 => q_2_port, IN2 => n8, QN => n10);
   U8 : NOR4X0 port map( IN1 => q_3_port, IN2 => n8, IN3 => n2, IN4 => n1, QN 
                           => n7);
   U9 : NOR2X0 port map( IN1 => q_0_port, IN2 => load, QN => n12);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_LWC_1.all;

entity xoodoo_round_ADDRESS_LEN128_ADDRESS_ENTRIES16_ADDRESS_ENTRIES_BITs4_1 is

   port( RAMA, RAMB : in std_logic_vector (127 downto 0);  perm_output : out 
         std_logic_vector (127 downto 0);  ADDRA, ADDRB : out std_logic_vector 
         (3 downto 0);  RNDCTR : in std_logic_vector (3 downto 0);  ins_counter
         : in std_logic_vector (4 downto 0));

end xoodoo_round_ADDRESS_LEN128_ADDRESS_ENTRIES16_ADDRESS_ENTRIES_BITs4_1;

architecture SYN_Behavioral of 
   xoodoo_round_ADDRESS_LEN128_ADDRESS_ENTRIES16_ADDRESS_ENTRIES_BITs4_1 is

   component NAND2X1
      port( IN1, IN2 : in std_logic;  QN : out std_logic);
   end component;
   
   component NAND3X0
      port( IN1, IN2, IN3 : in std_logic;  QN : out std_logic);
   end component;
   
   component OA22X1
      port( IN1, IN2, IN3, IN4 : in std_logic;  Q : out std_logic);
   end component;
   
   component OAI21X1
      port( IN1, IN2, IN3 : in std_logic;  QN : out std_logic);
   end component;
   
   component AO221X1
      port( IN1, IN2, IN3, IN4, IN5 : in std_logic;  Q : out std_logic);
   end component;
   
   component AO22X1
      port( IN1, IN2, IN3, IN4 : in std_logic;  Q : out std_logic);
   end component;
   
   component NOR2X0
      port( IN1, IN2 : in std_logic;  QN : out std_logic);
   end component;
   
   component NAND2X0
      port( IN1, IN2 : in std_logic;  QN : out std_logic);
   end component;
   
   component INVX0
      port( INP : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2X1
      port( IN1, IN2 : in std_logic;  Q : out std_logic);
   end component;
   
   component NBUFFX2
      port( INP : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2X4
      port( IN1, IN2 : in std_logic;  Q : out std_logic);
   end component;
   
   component XOR2X1
      port( IN1, IN2 : in std_logic;  Q : out std_logic);
   end component;
   
   component IBUFFX16
      port( INP : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2X2
      port( IN1, IN2 : in std_logic;  Q : out std_logic);
   end component;
   
   component DELLN1X2
      port( INP : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2X2
      port( IN1, IN2 : in std_logic;  Q : out std_logic);
   end component;
   
   component XNOR2X1
      port( IN1, IN2 : in std_logic;  Q : out std_logic);
   end component;
   
   component NAND4X0
      port( IN1, IN2, IN3, IN4 : in std_logic;  QN : out std_logic);
   end component;
   
   component AO21X1
      port( IN1, IN2, IN3 : in std_logic;  Q : out std_logic);
   end component;
   
   component AO222X1
      port( IN1, IN2, IN3, IN4, IN5, IN6 : in std_logic;  Q : out std_logic);
   end component;
   
   component OAI221X1
      port( IN1, IN2, IN3, IN4, IN5 : in std_logic;  QN : out std_logic);
   end component;
   
   component AND4X1
      port( IN1, IN2, IN3, IN4 : in std_logic;  Q : out std_logic);
   end component;
   
   component AND3X1
      port( IN1, IN2, IN3 : in std_logic;  Q : out std_logic);
   end component;
   
   component OA21X1
      port( IN1, IN2, IN3 : in std_logic;  Q : out std_logic);
   end component;
   
   component OR3X1
      port( IN1, IN2, IN3 : in std_logic;  Q : out std_logic);
   end component;
   
   component AOI22X1
      port( IN1, IN2, IN3, IN4 : in std_logic;  QN : out std_logic);
   end component;
   
   signal instruction_11_port, instruction_10_port, instruction_9_port, 
      instruction_8_port, addout_127_port, addout_126_port, addout_125_port, 
      addout_124_port, addout_123_port, addout_122_port, addout_121_port, 
      addout_120_port, addout_119_port, addout_118_port, addout_117_port, 
      addout_116_port, addout_115_port, addout_114_port, addout_113_port, 
      addout_112_port, addout_111_port, addout_110_port, addout_109_port, 
      addout_108_port, addout_107_port, addout_106_port, addout_105_port, 
      addout_104_port, addout_103_port, addout_102_port, addout_101_port, 
      addout_100_port, addout_99_port, addout_98_port, addout_97_port, 
      addout_96_port, addout_95_port, addout_94_port, addout_93_port, 
      addout_92_port, addout_91_port, addout_90_port, addout_89_port, 
      addout_88_port, addout_87_port, addout_86_port, addout_85_port, 
      addout_84_port, addout_83_port, addout_82_port, addout_81_port, 
      addout_80_port, addout_79_port, addout_78_port, addout_77_port, 
      addout_76_port, addout_75_port, addout_74_port, addout_73_port, 
      addout_72_port, addout_71_port, addout_70_port, addout_69_port, 
      addout_68_port, addout_67_port, addout_66_port, addout_65_port, 
      addout_64_port, addout_63_port, addout_62_port, addout_61_port, 
      addout_60_port, addout_59_port, addout_58_port, addout_57_port, 
      addout_56_port, addout_55_port, addout_54_port, addout_53_port, 
      addout_52_port, addout_51_port, addout_50_port, addout_49_port, 
      addout_48_port, addout_47_port, addout_46_port, addout_45_port, 
      addout_44_port, addout_43_port, addout_42_port, addout_41_port, 
      addout_40_port, addout_39_port, addout_38_port, addout_37_port, 
      addout_36_port, addout_35_port, addout_34_port, addout_33_port, 
      addout_32_port, addout_31_port, addout_30_port, addout_29_port, 
      addout_28_port, addout_27_port, addout_26_port, addout_25_port, 
      addout_24_port, addout_23_port, addout_22_port, addout_21_port, 
      addout_20_port, addout_19_port, addout_18_port, addout_17_port, 
      addout_16_port, addout_15_port, addout_14_port, addout_13_port, 
      addout_12_port, addout_11_port, addout_10_port, addout_9_port, 
      addout_8_port, addout_7_port, addout_6_port, addout_5_port, addout_4_port
      , addout_3_port, addout_2_port, addout_1_port, addout_0_port, 
      eshift_127_port, eshift_126_port, eshift_125_port, eshift_124_port, 
      eshift_123_port, eshift_122_port, eshift_121_port, eshift_120_port, 
      eshift_119_port, eshift_118_port, eshift_117_port, eshift_116_port, 
      eshift_115_port, eshift_114_port, eshift_113_port, eshift_112_port, 
      eshift_111_port, eshift_110_port, eshift_109_port, eshift_108_port, 
      eshift_107_port, eshift_106_port, eshift_105_port, eshift_104_port, 
      eshift_103_port, eshift_102_port, eshift_101_port, eshift_100_port, 
      eshift_99_port, eshift_98_port, eshift_97_port, eshift_96_port, 
      eshift_95_port, eshift_94_port, eshift_93_port, eshift_92_port, 
      eshift_91_port, eshift_90_port, eshift_89_port, eshift_88_port, 
      eshift_87_port, eshift_86_port, eshift_85_port, eshift_84_port, 
      eshift_83_port, eshift_82_port, eshift_81_port, eshift_80_port, 
      eshift_79_port, eshift_78_port, eshift_77_port, eshift_76_port, 
      eshift_75_port, eshift_74_port, eshift_73_port, eshift_72_port, 
      eshift_71_port, eshift_70_port, eshift_69_port, eshift_68_port, 
      eshift_67_port, eshift_66_port, eshift_65_port, eshift_64_port, 
      eshift_63_port, eshift_62_port, eshift_61_port, eshift_60_port, 
      eshift_59_port, eshift_58_port, eshift_57_port, eshift_56_port, 
      eshift_55_port, eshift_54_port, eshift_53_port, eshift_52_port, 
      eshift_51_port, eshift_50_port, eshift_49_port, eshift_48_port, 
      eshift_47_port, eshift_46_port, eshift_45_port, eshift_44_port, 
      eshift_43_port, eshift_42_port, eshift_41_port, eshift_40_port, 
      eshift_39_port, eshift_38_port, eshift_37_port, eshift_36_port, 
      eshift_35_port, eshift_34_port, eshift_33_port, eshift_32_port, 
      eshift_31_port, eshift_30_port, eshift_29_port, eshift_28_port, 
      eshift_27_port, eshift_26_port, eshift_25_port, eshift_24_port, 
      eshift_23_port, eshift_22_port, eshift_21_port, eshift_20_port, 
      eshift_19_port, eshift_18_port, eshift_17_port, eshift_16_port, 
      eshift_15_port, eshift_14_port, eshift_13_port, eshift_12_port, 
      eshift_11_port, eshift_10_port, eshift_9_port, eshift_8_port, 
      eshift_7_port, eshift_6_port, eshift_5_port, eshift_4_port, eshift_3_port
      , eshift_2_port, eshift_1_port, eshift_0_port, add_rnd_const_105_port, 
      add_rnd_const_104_port, add_rnd_const_103_port, add_rnd_const_102_port, 
      add_rnd_const_101_port, add_rnd_const_100_port, add_rnd_const_99_port, 
      add_rnd_const_98_port, add_rnd_const_97_port, andout_127_port, 
      andout_126_port, andout_125_port, andout_124_port, andout_123_port, 
      andout_122_port, andout_121_port, andout_120_port, andout_119_port, 
      andout_118_port, andout_117_port, andout_116_port, andout_115_port, 
      andout_114_port, andout_113_port, andout_112_port, andout_111_port, 
      andout_110_port, andout_109_port, andout_108_port, andout_107_port, 
      andout_106_port, andout_105_port, andout_104_port, andout_103_port, 
      andout_102_port, andout_101_port, andout_100_port, andout_99_port, 
      andout_98_port, andout_97_port, andout_96_port, andout_95_port, 
      andout_94_port, andout_93_port, andout_92_port, andout_91_port, 
      andout_90_port, andout_89_port, andout_88_port, andout_87_port, 
      andout_86_port, andout_85_port, andout_84_port, andout_83_port, 
      andout_82_port, andout_81_port, andout_80_port, andout_79_port, 
      andout_78_port, andout_77_port, andout_76_port, andout_75_port, 
      andout_74_port, andout_73_port, andout_72_port, andout_71_port, 
      andout_70_port, andout_69_port, andout_68_port, andout_67_port, 
      andout_66_port, andout_65_port, andout_64_port, andout_63_port, 
      andout_62_port, andout_61_port, andout_60_port, andout_59_port, 
      andout_58_port, andout_57_port, andout_56_port, andout_55_port, 
      andout_54_port, andout_53_port, andout_52_port, andout_51_port, 
      andout_50_port, andout_49_port, andout_48_port, andout_47_port, 
      andout_46_port, andout_45_port, andout_44_port, andout_43_port, 
      andout_42_port, andout_41_port, andout_40_port, andout_39_port, 
      andout_38_port, andout_37_port, andout_36_port, andout_35_port, 
      andout_34_port, andout_33_port, andout_32_port, andout_31_port, 
      andout_30_port, andout_29_port, andout_28_port, andout_27_port, 
      andout_26_port, andout_25_port, andout_24_port, andout_23_port, 
      andout_22_port, andout_21_port, andout_20_port, andout_19_port, 
      andout_18_port, andout_17_port, andout_16_port, andout_15_port, 
      andout_14_port, andout_13_port, andout_12_port, andout_11_port, 
      andout_10_port, andout_9_port, andout_8_port, andout_7_port, 
      andout_6_port, andout_5_port, andout_4_port, andout_3_port, andout_2_port
      , andout_1_port, andout_0_port, n145, n146, n147, n148, n149, n150, n151,
      n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, 
      n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, 
      n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, 
      n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, 
      n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, 
      n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31
      , n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, 
      n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60
      , n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, 
      n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89
      , n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, 
      n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, 
      n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, 
      n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, 
      n139, n140, n141, n142, n143, n144, n200, n201, n202, n203, n204, n205, 
      n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, 
      n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, 
      n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, 
      n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, 
      n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, 
      n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, 
      n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, 
      n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, 
      n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, 
      n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, 
      n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, 
      n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, 
      n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, 
      n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, 
      n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, 
      n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, 
      n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, 
      n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, 
      n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, 
      n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, 
      n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, 
      n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, 
      n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, 
      n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, 
      n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, 
      n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, 
      n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, 
      n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, 
      n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, 
      n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, 
      n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, 
      n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, 
      n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, 
      n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, 
      n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, 
      n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, 
      n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, 
      n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, 
      n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, 
      n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, 
      n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, 
      n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, 
      n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, 
      n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, 
      n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, 
      n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, 
      n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, 
      n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, 
      n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, 
      n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, 
      n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, 
      n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, 
      n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, 
      n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, 
      n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, 
      n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, 
      n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, 
      n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, 
      n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, 
      n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, 
      n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, 
      n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, 
      n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, 
      n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, 
      n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, 
      n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, 
      n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008
      , n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, 
      n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, 
      n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, 
      n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, 
      n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, 
      n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, 
      n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, 
      n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, 
      n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, 
      n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, 
      n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, 
      n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, 
      n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, 
      n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, 
      n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, 
      n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, 
      n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, 
      n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, 
      n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, 
      n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, 
      n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, 
      n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, 
      n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, 
      n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, 
      n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, 
      n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, 
      n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, 
      n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287 : std_logic
      ;

begin
   
   U178 : NAND3X0 port map( IN1 => n145, IN2 => n146, IN3 => n147, QN => 
                           instruction_9_port);
   U179 : NAND3X0 port map( IN1 => n149, IN2 => n150, IN3 => n151, QN => 
                           instruction_8_port);
   U180 : AOI22X1 port map( IN1 => n1272, IN2 => n152, IN3 => 
                           instruction_10_port, IN4 => ins_counter(0), QN => 
                           n151);
   U181 : OR3X1 port map( IN1 => n1143, IN2 => ins_counter(3), IN3 => n153, Q 
                           => n149);
   U182 : AO22X1 port map( IN1 => n1280, IN2 => n1272, IN3 => n154, IN4 => n152
                           , Q => instruction_11_port);
   U183 : XNOR2X1 port map( IN1 => n1203, IN2 => RAMB(36), Q => eshift_9_port);
   U184 : XNOR2X1 port map( IN1 => n1174, IN2 => RAMB(21), Q => eshift_99_port)
                           ;
   U185 : XNOR2X1 port map( IN1 => n1173, IN2 => RAMB(20), Q => eshift_98_port)
                           ;
   U186 : XNOR2X1 port map( IN1 => n1172, IN2 => RAMB(19), Q => eshift_97_port)
                           ;
   U187 : XNOR2X1 port map( IN1 => n1171, IN2 => RAMB(18), Q => eshift_96_port)
                           ;
   U188 : XNOR2X1 port map( IN1 => n1266, IN2 => RAMB(113), Q => eshift_95_port
                           );
   U189 : XNOR2X1 port map( IN1 => n1265, IN2 => RAMB(112), Q => eshift_94_port
                           );
   U190 : XNOR2X1 port map( IN1 => n1264, IN2 => RAMB(111), Q => eshift_93_port
                           );
   U191 : XNOR2X1 port map( IN1 => n1263, IN2 => RAMB(110), Q => eshift_92_port
                           );
   U192 : XNOR2X1 port map( IN1 => n1262, IN2 => RAMB(109), Q => eshift_91_port
                           );
   U193 : XNOR2X1 port map( IN1 => n1261, IN2 => RAMB(108), Q => eshift_90_port
                           );
   U194 : XNOR2X1 port map( IN1 => n1202, IN2 => RAMB(35), Q => eshift_8_port);
   U195 : XNOR2X1 port map( IN1 => n1260, IN2 => RAMB(107), Q => eshift_89_port
                           );
   U196 : XNOR2X1 port map( IN1 => n1259, IN2 => RAMB(106), Q => eshift_88_port
                           );
   U197 : XNOR2X1 port map( IN1 => n1258, IN2 => RAMB(105), Q => eshift_87_port
                           );
   U198 : XNOR2X1 port map( IN1 => n1257, IN2 => RAMB(104), Q => eshift_86_port
                           );
   U199 : XNOR2X1 port map( IN1 => n1256, IN2 => RAMB(103), Q => eshift_85_port
                           );
   U200 : XNOR2X1 port map( IN1 => n1255, IN2 => RAMB(102), Q => eshift_84_port
                           );
   U201 : XNOR2X1 port map( IN1 => n1254, IN2 => RAMB(101), Q => eshift_83_port
                           );
   U202 : XNOR2X1 port map( IN1 => n1253, IN2 => RAMB(100), Q => eshift_82_port
                           );
   U203 : XNOR2X1 port map( IN1 => n1243, IN2 => RAMB(108), Q => eshift_81_port
                           );
   U204 : XNOR2X1 port map( IN1 => n1242, IN2 => RAMB(107), Q => eshift_80_port
                           );
   U205 : XNOR2X1 port map( IN1 => n1201, IN2 => RAMB(34), Q => eshift_7_port);
   U206 : XNOR2X1 port map( IN1 => n1241, IN2 => RAMB(106), Q => eshift_79_port
                           );
   U207 : XNOR2X1 port map( IN1 => n1240, IN2 => RAMB(105), Q => eshift_78_port
                           );
   U208 : XNOR2X1 port map( IN1 => n1271, IN2 => RAMB(104), Q => eshift_77_port
                           );
   U209 : XNOR2X1 port map( IN1 => n1270, IN2 => RAMB(103), Q => eshift_76_port
                           );
   U210 : XNOR2X1 port map( IN1 => n1269, IN2 => RAMB(102), Q => eshift_75_port
                           );
   U211 : XNOR2X1 port map( IN1 => n1268, IN2 => RAMB(101), Q => eshift_74_port
                           );
   U212 : XNOR2X1 port map( IN1 => n1267, IN2 => RAMB(100), Q => eshift_73_port
                           );
   U213 : XNOR2X1 port map( IN1 => n1243, IN2 => RAMB(122), Q => eshift_72_port
                           );
   U214 : XNOR2X1 port map( IN1 => n1242, IN2 => RAMB(121), Q => eshift_71_port
                           );
   U215 : XNOR2X1 port map( IN1 => n1241, IN2 => RAMB(120), Q => eshift_70_port
                           );
   U216 : XNOR2X1 port map( IN1 => n1200, IN2 => RAMB(33), Q => eshift_6_port);
   U217 : XNOR2X1 port map( IN1 => n1240, IN2 => RAMB(119), Q => eshift_69_port
                           );
   U218 : XNOR2X1 port map( IN1 => n1271, IN2 => RAMB(118), Q => eshift_68_port
                           );
   U219 : XNOR2X1 port map( IN1 => n1270, IN2 => RAMB(117), Q => eshift_67_port
                           );
   U220 : XNOR2X1 port map( IN1 => n1269, IN2 => RAMB(116), Q => eshift_66_port
                           );
   U221 : XNOR2X1 port map( IN1 => n1268, IN2 => RAMB(115), Q => eshift_65_port
                           );
   U222 : XNOR2X1 port map( IN1 => n1267, IN2 => RAMB(114), Q => eshift_64_port
                           );
   U223 : XNOR2X1 port map( IN1 => n1234, IN2 => RAMB(81), Q => eshift_63_port)
                           ;
   U224 : XNOR2X1 port map( IN1 => n1233, IN2 => RAMB(80), Q => eshift_62_port)
                           ;
   U225 : XNOR2X1 port map( IN1 => n1232, IN2 => RAMB(79), Q => eshift_61_port)
                           ;
   U226 : XNOR2X1 port map( IN1 => n1231, IN2 => RAMB(78), Q => eshift_60_port)
                           ;
   U227 : XNOR2X1 port map( IN1 => n1199, IN2 => RAMB(32), Q => eshift_5_port);
   U228 : XNOR2X1 port map( IN1 => n1230, IN2 => RAMB(77), Q => eshift_59_port)
                           ;
   U229 : XNOR2X1 port map( IN1 => n1229, IN2 => RAMB(76), Q => eshift_58_port)
                           ;
   U230 : XNOR2X1 port map( IN1 => n1228, IN2 => RAMB(75), Q => eshift_57_port)
                           ;
   U231 : XNOR2X1 port map( IN1 => n1227, IN2 => RAMB(74), Q => eshift_56_port)
                           ;
   U232 : XNOR2X1 port map( IN1 => n1226, IN2 => RAMB(73), Q => eshift_55_port)
                           ;
   U233 : XNOR2X1 port map( IN1 => n1225, IN2 => RAMB(72), Q => eshift_54_port)
                           ;
   U234 : XNOR2X1 port map( IN1 => n1224, IN2 => RAMB(71), Q => eshift_53_port)
                           ;
   U235 : XNOR2X1 port map( IN1 => n1223, IN2 => RAMB(70), Q => eshift_52_port)
                           ;
   U236 : XNOR2X1 port map( IN1 => n1222, IN2 => RAMB(69), Q => eshift_51_port)
                           ;
   U237 : XNOR2X1 port map( IN1 => n1221, IN2 => RAMB(68), Q => eshift_50_port)
                           ;
   U238 : XNOR2X1 port map( IN1 => n1207, IN2 => RAMB(54), Q => eshift_4_port);
   U239 : XNOR2X1 port map( IN1 => n1220, IN2 => RAMB(67), Q => eshift_49_port)
                           ;
   U240 : XNOR2X1 port map( IN1 => n1219, IN2 => RAMB(66), Q => eshift_48_port)
                           ;
   U241 : XNOR2X1 port map( IN1 => n1218, IN2 => RAMB(65), Q => eshift_47_port)
                           ;
   U242 : XNOR2X1 port map( IN1 => n1217, IN2 => RAMB(64), Q => eshift_46_port)
                           ;
   U243 : XNOR2X1 port map( IN1 => n1239, IN2 => RAMB(72), Q => eshift_45_port)
                           ;
   U244 : XNOR2X1 port map( IN1 => n1238, IN2 => RAMB(71), Q => eshift_44_port)
                           ;
   U245 : XNOR2X1 port map( IN1 => n1237, IN2 => RAMB(70), Q => eshift_43_port)
                           ;
   U246 : XNOR2X1 port map( IN1 => n1236, IN2 => RAMB(69), Q => eshift_42_port)
                           ;
   U247 : XNOR2X1 port map( IN1 => n1235, IN2 => RAMB(68), Q => eshift_41_port)
                           ;
   U248 : XNOR2X1 port map( IN1 => n1234, IN2 => RAMB(67), Q => eshift_40_port)
                           ;
   U249 : XNOR2X1 port map( IN1 => n1206, IN2 => RAMB(53), Q => eshift_3_port);
   U250 : XNOR2X1 port map( IN1 => n1233, IN2 => RAMB(66), Q => eshift_39_port)
                           ;
   U251 : XNOR2X1 port map( IN1 => n1232, IN2 => RAMB(65), Q => eshift_38_port)
                           ;
   U252 : XNOR2X1 port map( IN1 => n1231, IN2 => RAMB(64), Q => eshift_37_port)
                           ;
   U253 : XNOR2X1 port map( IN1 => n1239, IN2 => RAMB(86), Q => eshift_36_port)
                           ;
   U254 : XNOR2X1 port map( IN1 => n1238, IN2 => RAMB(85), Q => eshift_35_port)
                           ;
   U255 : XNOR2X1 port map( IN1 => n1237, IN2 => RAMB(84), Q => eshift_34_port)
                           ;
   U256 : XNOR2X1 port map( IN1 => n1236, IN2 => RAMB(83), Q => eshift_33_port)
                           ;
   U257 : XNOR2X1 port map( IN1 => n1235, IN2 => RAMB(82), Q => eshift_32_port)
                           ;
   U258 : XNOR2X1 port map( IN1 => n1202, IN2 => RAMB(49), Q => eshift_31_port)
                           ;
   U259 : XNOR2X1 port map( IN1 => n1201, IN2 => RAMB(48), Q => eshift_30_port)
                           ;
   U260 : XNOR2X1 port map( IN1 => n1205, IN2 => RAMB(52), Q => eshift_2_port);
   U261 : XNOR2X1 port map( IN1 => n1200, IN2 => RAMB(47), Q => eshift_29_port)
                           ;
   U262 : XNOR2X1 port map( IN1 => n1199, IN2 => RAMB(46), Q => eshift_28_port)
                           ;
   U263 : XNOR2X1 port map( IN1 => n1198, IN2 => RAMB(45), Q => eshift_27_port)
                           ;
   U264 : XNOR2X1 port map( IN1 => n1197, IN2 => RAMB(44), Q => eshift_26_port)
                           ;
   U265 : XNOR2X1 port map( IN1 => n1196, IN2 => RAMB(43), Q => eshift_25_port)
                           ;
   U266 : XNOR2X1 port map( IN1 => n1195, IN2 => RAMB(42), Q => eshift_24_port)
                           ;
   U267 : XNOR2X1 port map( IN1 => n1194, IN2 => RAMB(41), Q => eshift_23_port)
                           ;
   U268 : XNOR2X1 port map( IN1 => n1193, IN2 => RAMB(40), Q => eshift_22_port)
                           ;
   U269 : XNOR2X1 port map( IN1 => n1192, IN2 => RAMB(39), Q => eshift_21_port)
                           ;
   U270 : XNOR2X1 port map( IN1 => n1191, IN2 => RAMB(38), Q => eshift_20_port)
                           ;
   U271 : XNOR2X1 port map( IN1 => n1204, IN2 => RAMB(51), Q => eshift_1_port);
   U272 : XNOR2X1 port map( IN1 => n1190, IN2 => RAMB(37), Q => eshift_19_port)
                           ;
   U273 : XNOR2X1 port map( IN1 => n1189, IN2 => n17, Q => eshift_18_port);
   U274 : XNOR2X1 port map( IN1 => n1188, IN2 => RAMB(35), Q => eshift_17_port)
                           ;
   U275 : XNOR2X1 port map( IN1 => n1187, IN2 => RAMB(34), Q => eshift_16_port)
                           ;
   U276 : XNOR2X1 port map( IN1 => n1186, IN2 => RAMB(33), Q => eshift_15_port)
                           ;
   U277 : XNOR2X1 port map( IN1 => n1185, IN2 => RAMB(32), Q => eshift_14_port)
                           ;
   U278 : XNOR2X1 port map( IN1 => n1207, IN2 => RAMB(40), Q => eshift_13_port)
                           ;
   U279 : XNOR2X1 port map( IN1 => n1206, IN2 => n16, Q => eshift_12_port);
   U280 : XNOR2X1 port map( IN1 => n1170, IN2 => RAMB(17), Q => eshift_127_port
                           );
   U281 : XNOR2X1 port map( IN1 => n1169, IN2 => RAMB(16), Q => eshift_126_port
                           );
   U282 : XNOR2X1 port map( IN1 => n1168, IN2 => RAMB(15), Q => eshift_125_port
                           );
   U283 : XNOR2X1 port map( IN1 => n1167, IN2 => RAMB(14), Q => eshift_124_port
                           );
   U284 : XNOR2X1 port map( IN1 => n1166, IN2 => RAMB(13), Q => eshift_123_port
                           );
   U285 : XNOR2X1 port map( IN1 => n1165, IN2 => RAMB(12), Q => eshift_122_port
                           );
   U286 : XNOR2X1 port map( IN1 => n1164, IN2 => RAMB(11), Q => eshift_121_port
                           );
   U287 : XNOR2X1 port map( IN1 => n1163, IN2 => RAMB(10), Q => eshift_120_port
                           );
   U288 : XNOR2X1 port map( IN1 => n1205, IN2 => RAMB(38), Q => eshift_11_port)
                           ;
   U289 : XNOR2X1 port map( IN1 => n1153, IN2 => RAMB(18), Q => eshift_119_port
                           );
   U290 : XNOR2X1 port map( IN1 => n1152, IN2 => RAMB(17), Q => eshift_118_port
                           );
   U291 : XNOR2X1 port map( IN1 => n1151, IN2 => RAMB(16), Q => eshift_117_port
                           );
   U292 : XNOR2X1 port map( IN1 => n1150, IN2 => RAMB(15), Q => eshift_116_port
                           );
   U293 : XNOR2X1 port map( IN1 => n1149, IN2 => RAMB(14), Q => eshift_115_port
                           );
   U294 : XNOR2X1 port map( IN1 => n1148, IN2 => RAMB(13), Q => eshift_114_port
                           );
   U295 : XNOR2X1 port map( IN1 => n1147, IN2 => RAMB(12), Q => eshift_113_port
                           );
   U296 : XNOR2X1 port map( IN1 => n1146, IN2 => RAMB(11), Q => eshift_112_port
                           );
   U297 : XNOR2X1 port map( IN1 => n1145, IN2 => RAMB(10), Q => eshift_111_port
                           );
   U298 : XNOR2X1 port map( IN1 => n1153, IN2 => RAMB(0), Q => eshift_110_port)
                           ;
   U299 : XNOR2X1 port map( IN1 => n1204, IN2 => RAMB(37), Q => eshift_10_port)
                           ;
   U300 : XNOR2X1 port map( IN1 => n1152, IN2 => RAMB(31), Q => eshift_109_port
                           );
   U301 : XNOR2X1 port map( IN1 => n1151, IN2 => RAMB(30), Q => eshift_108_port
                           );
   U302 : XNOR2X1 port map( IN1 => n1150, IN2 => RAMB(29), Q => eshift_107_port
                           );
   U303 : XNOR2X1 port map( IN1 => n1149, IN2 => RAMB(28), Q => eshift_106_port
                           );
   U304 : XNOR2X1 port map( IN1 => n1148, IN2 => RAMB(27), Q => eshift_105_port
                           );
   U305 : XNOR2X1 port map( IN1 => n1147, IN2 => RAMB(26), Q => eshift_104_port
                           );
   U306 : XNOR2X1 port map( IN1 => n1146, IN2 => RAMB(25), Q => eshift_103_port
                           );
   U307 : XNOR2X1 port map( IN1 => n1168, IN2 => RAMB(1), Q => eshift_102_port)
                           ;
   U308 : XNOR2X1 port map( IN1 => n1167, IN2 => RAMB(0), Q => eshift_101_port)
                           ;
   U309 : XNOR2X1 port map( IN1 => n1175, IN2 => RAMB(22), Q => eshift_100_port
                           );
   U310 : XNOR2X1 port map( IN1 => n1203, IN2 => RAMB(50), Q => eshift_0_port);
   U316 : AND2X1 port map( IN1 => RAMB(95), IN2 => n212, Q => andout_95_port);
   U319 : AND2X1 port map( IN1 => RAMB(92), IN2 => n218, Q => andout_92_port);
   U324 : AND2X1 port map( IN1 => RAMB(88), IN2 => n217, Q => andout_88_port);
   U339 : AND2X1 port map( IN1 => RAMB(74), IN2 => n139, Q => andout_74_port);
   U348 : AND2X1 port map( IN1 => RAMB(66), IN2 => n223, Q => andout_66_port);
   U384 : AND2X1 port map( IN1 => RAMB(33), IN2 => n141, Q => andout_33_port);
   U388 : AND2X1 port map( IN1 => RAMB(2), IN2 => n208, Q => andout_2_port);
   U392 : AND2X1 port map( IN1 => RAMB(26), IN2 => n205, Q => andout_26_port);
   U396 : AND2X1 port map( IN1 => RAMB(22), IN2 => n210, Q => andout_22_port);
   U397 : AND2X1 port map( IN1 => RAMB(21), IN2 => n201, Q => andout_21_port);
   U412 : AND2X1 port map( IN1 => RAMB(123), IN2 => n222, Q => andout_123_port)
                           ;
   U421 : AND2X1 port map( IN1 => RAMB(115), IN2 => n26, Q => andout_115_port);
   U429 : AND2X1 port map( IN1 => RAMB(108), IN2 => n213, Q => andout_108_port)
                           ;
   U439 : XNOR2X1 port map( IN1 => n1153, IN2 => n92, Q => addout_9_port);
   U440 : XNOR2X1 port map( IN1 => n1243, IN2 => n34, Q => addout_99_port);
   U443 : XNOR2X1 port map( IN1 => n1240, IN2 => n114, Q => addout_96_port);
   U445 : XNOR2X1 port map( IN1 => n1238, IN2 => n113, Q => addout_94_port);
   U448 : XNOR2X1 port map( IN1 => n1235, IN2 => n71, Q => addout_91_port);
   U449 : XNOR2X1 port map( IN1 => n1234, IN2 => n123, Q => addout_90_port);
   U450 : XNOR2X1 port map( IN1 => n1152, IN2 => n102, Q => addout_8_port);
   U451 : XNOR2X1 port map( IN1 => n1233, IN2 => n66, Q => addout_89_port);
   U453 : XNOR2X1 port map( IN1 => n1231, IN2 => n77, Q => addout_87_port);
   U454 : XNOR2X1 port map( IN1 => n1230, IN2 => n95, Q => addout_86_port);
   U457 : XNOR2X1 port map( IN1 => n1227, IN2 => n63, Q => addout_83_port);
   U458 : XNOR2X1 port map( IN1 => n105, IN2 => n1226, Q => addout_82_port);
   U459 : XNOR2X1 port map( IN1 => n118, IN2 => n1225, Q => addout_81_port);
   U460 : XNOR2X1 port map( IN1 => n1224, IN2 => n56, Q => addout_80_port);
   U461 : XNOR2X1 port map( IN1 => n111, IN2 => n1151, Q => addout_7_port);
   U462 : XNOR2X1 port map( IN1 => n1223, IN2 => n115, Q => addout_79_port);
   U463 : XNOR2X1 port map( IN1 => n1222, IN2 => n107, Q => addout_78_port);
   U464 : XNOR2X1 port map( IN1 => n62, IN2 => n1221, Q => addout_77_port);
   U465 : XNOR2X1 port map( IN1 => n137, IN2 => n1220, Q => addout_76_port);
   U466 : XNOR2X1 port map( IN1 => n42, IN2 => n1219, Q => addout_75_port);
   U467 : XNOR2X1 port map( IN1 => n1218, IN2 => n27, Q => addout_74_port);
   U468 : XNOR2X1 port map( IN1 => n1217, IN2 => n110, Q => addout_73_port);
   U469 : XNOR2X1 port map( IN1 => n1216, IN2 => n128, Q => addout_72_port);
   U471 : XNOR2X1 port map( IN1 => n58, IN2 => n1214, Q => addout_70_port);
   U472 : XNOR2X1 port map( IN1 => n135, IN2 => n1150, Q => addout_6_port);
   U473 : XNOR2X1 port map( IN1 => n109, IN2 => n1213, Q => addout_69_port);
   U475 : XNOR2X1 port map( IN1 => n79, IN2 => n1211, Q => addout_67_port);
   U477 : XNOR2X1 port map( IN1 => n49, IN2 => n1209, Q => addout_65_port);
   U478 : XNOR2X1 port map( IN1 => n121, IN2 => n1208, Q => addout_64_port);
   U479 : XNOR2X1 port map( IN1 => n1207, IN2 => n78, Q => addout_63_port);
   U480 : XNOR2X1 port map( IN1 => n52, IN2 => n1206, Q => addout_62_port);
   U481 : XNOR2X1 port map( IN1 => n1205, IN2 => n100, Q => addout_61_port);
   U482 : XNOR2X1 port map( IN1 => n1204, IN2 => n81, Q => addout_60_port);
   U484 : XNOR2X1 port map( IN1 => n1203, IN2 => n53, Q => addout_59_port);
   U485 : XNOR2X1 port map( IN1 => n124, IN2 => n1202, Q => addout_58_port);
   U487 : XNOR2X1 port map( IN1 => n1200, IN2 => n136, Q => addout_56_port);
   U488 : XNOR2X1 port map( IN1 => n1199, IN2 => n69, Q => addout_55_port);
   U490 : XNOR2X1 port map( IN1 => n131, IN2 => n1197, Q => addout_53_port);
   U491 : XNOR2X1 port map( IN1 => n31, IN2 => n1196, Q => addout_52_port);
   U492 : XNOR2X1 port map( IN1 => n1195, IN2 => n133, Q => addout_51_port);
   U493 : XNOR2X1 port map( IN1 => n1194, IN2 => n116, Q => addout_50_port);
   U494 : XNOR2X1 port map( IN1 => n89, IN2 => n1148, Q => addout_4_port);
   U497 : XNOR2X1 port map( IN1 => n1191, IN2 => n134, Q => addout_47_port);
   U498 : XNOR2X1 port map( IN1 => n85, IN2 => n1190, Q => addout_46_port);
   U499 : XNOR2X1 port map( IN1 => n1189, IN2 => n67, Q => addout_45_port);
   U501 : XNOR2X1 port map( IN1 => n40, IN2 => n1187, Q => addout_43_port);
   U502 : XNOR2X1 port map( IN1 => n82, IN2 => n1186, Q => addout_42_port);
   U503 : XNOR2X1 port map( IN1 => n61, IN2 => n1185, Q => addout_41_port);
   U504 : XNOR2X1 port map( IN1 => n1184, IN2 => n74, Q => addout_40_port);
   U507 : XNOR2X1 port map( IN1 => n120, IN2 => n1182, Q => addout_38_port);
   U508 : XNOR2X1 port map( IN1 => n1181, IN2 => n48, Q => addout_37_port);
   U511 : XNOR2X1 port map( IN1 => n108, IN2 => n1178, Q => addout_34_port);
   U514 : XNOR2X1 port map( IN1 => n1175, IN2 => n98, Q => addout_31_port);
   U515 : XNOR2X1 port map( IN1 => n1174, IN2 => n37, Q => addout_30_port);
   U517 : XNOR2X1 port map( IN1 => n1173, IN2 => n126, Q => addout_29_port);
   U518 : XNOR2X1 port map( IN1 => n1172, IN2 => n119, Q => addout_28_port);
   U519 : XNOR2X1 port map( IN1 => n1171, IN2 => n68, Q => addout_27_port);
   U521 : XNOR2X1 port map( IN1 => n1169, IN2 => n73, Q => addout_25_port);
   U522 : XNOR2X1 port map( IN1 => n1168, IN2 => n36, Q => addout_24_port);
   U525 : XNOR2X1 port map( IN1 => n1165, IN2 => n35, Q => addout_21_port);
   U526 : XNOR2X1 port map( IN1 => n1164, IN2 => n132, Q => addout_20_port);
   U528 : XNOR2X1 port map( IN1 => n1163, IN2 => n72, Q => addout_19_port);
   U529 : XNOR2X1 port map( IN1 => n1162, IN2 => n55, Q => addout_18_port);
   U530 : XNOR2X1 port map( IN1 => n122, IN2 => n1161, Q => addout_17_port);
   U531 : XNOR2X1 port map( IN1 => n1160, IN2 => n117, Q => addout_16_port);
   U532 : XNOR2X1 port map( IN1 => n101, IN2 => n1159, Q => addout_15_port);
   U533 : XNOR2X1 port map( IN1 => n125, IN2 => n1158, Q => addout_14_port);
   U534 : XNOR2X1 port map( IN1 => n1157, IN2 => n127, Q => addout_13_port);
   U535 : XNOR2X1 port map( IN1 => n1156, IN2 => n75, Q => addout_12_port);
   U536 : XNOR2X1 port map( IN1 => n1271, IN2 => n28, Q => addout_127_port);
   U538 : XNOR2X1 port map( IN1 => n1269, IN2 => n76, Q => addout_125_port);
   U539 : XNOR2X1 port map( IN1 => n1268, IN2 => n50, Q => addout_124_port);
   U541 : XNOR2X1 port map( IN1 => n1266, IN2 => n96, Q => addout_122_port);
   U543 : XNOR2X1 port map( IN1 => n1264, IN2 => n2, Q => addout_120_port);
   U544 : XNOR2X1 port map( IN1 => n97, IN2 => n1155, Q => addout_11_port);
   U545 : XNOR2X1 port map( IN1 => n47, IN2 => n1263, Q => addout_119_port);
   U546 : XNOR2X1 port map( IN1 => n1262, IN2 => n80, Q => addout_118_port);
   U549 : XNOR2X1 port map( IN1 => n1259, IN2 => n26, Q => addout_115_port);
   U550 : XNOR2X1 port map( IN1 => n1258, IN2 => n103, Q => addout_114_port);
   U551 : XNOR2X1 port map( IN1 => n1257, IN2 => n57, Q => addout_113_port);
   U553 : XNOR2X1 port map( IN1 => n41, IN2 => n1255, Q => addout_111_port);
   U555 : XNOR2X1 port map( IN1 => n93, IN2 => n1154, Q => addout_10_port);
   U558 : XNOR2X1 port map( IN1 => n87, IN2 => n1251, Q => addout_107_port);
   U559 : XNOR2X1 port map( IN1 => n1250, IN2 => n106, Q => addout_106_port);
   U561 : XNOR2X1 port map( IN1 => n1248, IN2 => n144, Q => addout_104_port);
   U563 : XNOR2X1 port map( IN1 => n88, IN2 => n1246, Q => addout_102_port);
   U564 : XNOR2X1 port map( IN1 => n1245, IN2 => n94, Q => addout_101_port);
   U567 : XOR2X1 port map( IN1 => n156, IN2 => n34, Q => add_rnd_const_99_port)
                           ;
   U568 : NAND3X0 port map( IN1 => n157, IN2 => n158, IN3 => n159, QN => n156);
   U572 : OA21X1 port map( IN1 => RNDCTR(1), IN2 => n164, IN3 => n165, Q => 
                           n163);
   U573 : XOR2X1 port map( IN1 => n166, IN2 => n203, Q => 
                           add_rnd_const_104_port);
   U574 : NAND3X0 port map( IN1 => n164, IN2 => n165, IN3 => n167, QN => n166);
   U575 : NAND3X0 port map( IN1 => n1284, IN2 => n1286, IN3 => RNDCTR(2), QN =>
                           n167);
   U576 : XOR2X1 port map( IN1 => n168, IN2 => n86, Q => add_rnd_const_103_port
                           );
   U577 : NAND4X0 port map( IN1 => n164, IN2 => n169, IN3 => n170, IN4 => n165,
                           QN => n168);
   U578 : XOR2X1 port map( IN1 => n171, IN2 => n88, Q => add_rnd_const_102_port
                           );
   U579 : NAND3X0 port map( IN1 => n172, IN2 => n165, IN3 => n173, QN => n171);
   U580 : NAND3X0 port map( IN1 => n174, IN2 => n1284, IN3 => RNDCTR(1), QN => 
                           n165);
   U581 : XOR2X1 port map( IN1 => n175, IN2 => n94, Q => add_rnd_const_101_port
                           );
   U582 : NAND4X0 port map( IN1 => n169, IN2 => n157, IN3 => n1285, IN4 => n176
                           , QN => n175);
   U583 : OA22X1 port map( IN1 => n1286, IN2 => n164, IN3 => RNDCTR(0), IN4 => 
                           n1287, Q => n176);
   U584 : XOR2X1 port map( IN1 => n178, IN2 => n143, Q => 
                           add_rnd_const_100_port);
   U585 : NAND3X0 port map( IN1 => n1283, IN2 => n162, IN3 => n173, QN => n178)
                           ;
   U586 : AND3X1 port map( IN1 => n170, IN2 => n158, IN3 => n169, Q => n173);
   U587 : NAND3X0 port map( IN1 => n1284, IN2 => n1286, IN3 => n174, QN => n158
                           );
   U588 : NAND3X0 port map( IN1 => RNDCTR(0), IN2 => n174, IN3 => RNDCTR(1), QN
                           => n170);
   U589 : NAND3X0 port map( IN1 => RNDCTR(1), IN2 => RNDCTR(0), IN3 => 
                           RNDCTR(3), QN => n162);
   U590 : AND4X1 port map( IN1 => n1278, IN2 => ins_counter(3), IN3 => 
                           ins_counter(4), IN4 => n179, Q => ADDRB(3));
   U591 : NAND3X0 port map( IN1 => n180, IN2 => n181, IN3 => n182, QN => 
                           ADDRB(2));
   U592 : OA22X1 port map( IN1 => n148, IN2 => n150, IN3 => n1142, IN4 => n183,
                           Q => n182);
   U593 : AO221X1 port map( IN1 => n1280, IN2 => n153, IN3 => n184, IN4 => 
                           n1278, IN5 => n185, Q => ADDRB(1));
   U594 : OAI21X1 port map( IN1 => n145, IN2 => n155, IN3 => n181, QN => n185);
   U595 : AO222X1 port map( IN1 => n186, IN2 => n1274, IN3 => n187, IN4 => 
                           ins_counter(1), IN5 => instruction_10_port, IN6 => 
                           n153, Q => n184);
   U596 : NAND3X0 port map( IN1 => n189, IN2 => n183, IN3 => n190, QN => 
                           ADDRB(0));
   U597 : OA22X1 port map( IN1 => n1143, IN2 => n191, IN3 => n1274, IN4 => n181
                           , Q => n190);
   U598 : NAND3X0 port map( IN1 => ins_counter(3), IN2 => n1278, IN3 => n186, 
                           QN => n181);
   U599 : OA22X1 port map( IN1 => n1274, IN2 => n192, IN3 => ins_counter(0), 
                           IN4 => n193, Q => n191);
   U600 : NAND3X0 port map( IN1 => n1142, IN2 => n1282, IN3 => n148, QN => n189
                           );
   U601 : OAI221X1 port map( IN1 => n188, IN2 => n153, IN3 => n194, IN4 => 
                           n1273, IN5 => n145, QN => ADDRA(2));
   U602 : AO222X1 port map( IN1 => n195, IN2 => n1278, IN3 => n196, IN4 => 
                           n1275, IN5 => n179, IN6 => n1281, Q => ADDRA(1));
   U603 : AO21X1 port map( IN1 => n1276, IN2 => n1274, IN3 => n1277, Q => n195)
                           ;
   U604 : NAND4X0 port map( IN1 => n180, IN2 => n146, IN3 => n197, IN4 => n198,
                           QN => ADDRA(0));
   U605 : OA22X1 port map( IN1 => ins_counter(0), IN2 => n194, IN3 => n1278, 
                           IN4 => n183, Q => n198);
   U606 : AO221X1 port map( IN1 => n187, IN2 => n1275, IN3 => n152, IN4 => 
                           n1278, IN5 => n1279, Q => n199);
   U607 : NAND3X0 port map( IN1 => ins_counter(0), IN2 => n1278, IN3 => n186, 
                           QN => n180);
   U3 : NBUFFX2 port map( INP => RAMA(124), Z => n50);
   U4 : XOR2X1 port map( IN1 => RAMB(109), IN2 => n104, Q => addout_109_port);
   U5 : AND2X4 port map( IN1 => RAMB(109), IN2 => n104, Q => andout_109_port);
   U6 : NBUFFX2 port map( INP => RAMA(80), Z => n56);
   U7 : INVX0 port map( INP => n20, ZN => n1);
   U8 : INVX0 port map( INP => RAMA(48), ZN => n20);
   U9 : NBUFFX2 port map( INP => RAMA(24), Z => n36);
   U10 : NAND2X0 port map( IN1 => n365, IN2 => n6, QN => perm_output(105));
   U11 : XOR2X1 port map( IN1 => n1261, IN2 => n45, Q => addout_117_port);
   U12 : INVX0 port map( INP => RAMA(88), ZN => n216);
   U13 : NBUFFX2 port map( INP => RAMA(122), Z => n96);
   U14 : NBUFFX2 port map( INP => RAMA(106), Z => n106);
   U15 : NBUFFX2 port map( INP => RAMA(40), Z => n74);
   U16 : NBUFFX2 port map( INP => RAMA(16), Z => n117);
   U17 : NBUFFX2 port map( INP => RAMA(72), Z => n128);
   U18 : NBUFFX2 port map( INP => RAMA(61), Z => n100);
   U19 : INVX0 port map( INP => RAMA(21), ZN => n200);
   U20 : NBUFFX2 port map( INP => RAMA(73), Z => n110);
   U21 : NBUFFX2 port map( INP => RAMA(25), Z => n73);
   U22 : AND2X4 port map( IN1 => RAMB(126), IN2 => RAMA(126), Q => 
                           andout_126_port);
   U23 : NBUFFX2 port map( INP => RAMA(120), Z => n2);
   U24 : INVX0 port map( INP => RAMA(105), ZN => n3);
   U25 : INVX0 port map( INP => n3, ZN => n4);
   U26 : NBUFFX2 port map( INP => RAMA(56), Z => n136);
   U27 : XOR2X2 port map( IN1 => n7, IN2 => n1256, Q => addout_112_port);
   U28 : NAND2X1 port map( IN1 => n364, IN2 => n1128, QN => n5);
   U29 : INVX0 port map( INP => n5, ZN => n6);
   U30 : INVX0 port map( INP => RAMA(94), ZN => n112);
   U31 : NBUFFX2 port map( INP => RAMA(8), Z => n102);
   U32 : NBUFFX2 port map( INP => RAMA(10), Z => n93);
   U33 : NBUFFX2 port map( INP => RAMA(109), Z => n104);
   U34 : INVX0 port map( INP => RAMA(89), ZN => n65);
   U35 : NBUFFX2 port map( INP => RAMA(42), Z => n82);
   U36 : NBUFFX2 port map( INP => RAMA(30), Z => n37);
   U37 : XOR2X1 port map( IN1 => n206, IN2 => n1201, Q => addout_57_port);
   U38 : INVX0 port map( INP => RAMA(112), ZN => n7);
   U39 : INVX0 port map( INP => n7, ZN => n8);
   U40 : NBUFFX2 port map( INP => RAMA(13), Z => n127);
   U41 : NBUFFX2 port map( INP => RAMA(45), Z => n67);
   U42 : XNOR2X1 port map( IN1 => n19, IN2 => n1215, Q => addout_71_port);
   U43 : AND2X1 port map( IN1 => n952, IN2 => n1005, Q => n9);
   U44 : AND2X1 port map( IN1 => n244, IN2 => n1129, Q => n10);
   U45 : AND2X1 port map( IN1 => n466, IN2 => n1126, Q => n11);
   U46 : AND2X1 port map( IN1 => n652, IN2 => n1124, Q => n12);
   U47 : AND2X1 port map( IN1 => n544, IN2 => n1125, Q => n13);
   U48 : AND2X1 port map( IN1 => n232, IN2 => n1129, Q => n14);
   U49 : AND2X1 port map( IN1 => n862, IN2 => n1123, Q => n15);
   U50 : NBUFFX2 port map( INP => RAMA(37), Z => n48);
   U51 : NBUFFX2 port map( INP => RAMA(43), Z => n40);
   U52 : NBUFFX2 port map( INP => RAMA(52), Z => n31);
   U53 : NBUFFX2 port map( INP => RAMA(99), Z => n34);
   U54 : XOR2X2 port map( IN1 => n24, IN2 => n1241, Q => addout_97_port);
   U55 : INVX0 port map( INP => n1183, ZN => n16);
   U56 : INVX0 port map( INP => n1180, ZN => n17);
   U57 : XOR2X1 port map( IN1 => n16, IN2 => n64, Q => addout_39_port);
   U58 : XOR2X1 port map( IN1 => RAMB(5), IN2 => n60, Q => addout_5_port);
   U59 : XOR2X1 port map( IN1 => n17, IN2 => n129, Q => addout_36_port);
   U60 : XOR2X2 port map( IN1 => n142, IN2 => n1244, Q => addout_100_port);
   U61 : XNOR2X1 port map( IN1 => n25, IN2 => n162, Q => add_rnd_const_97_port)
                           ;
   U62 : AND2X1 port map( IN1 => RAMB(103), IN2 => n86, Q => andout_103_port);
   U63 : XOR2X2 port map( IN1 => n22, IN2 => n1242, Q => addout_98_port);
   U64 : XOR2X2 port map( IN1 => RAMB(66), IN2 => n223, Q => addout_66_port);
   U65 : NBUFFX2 port map( INP => RAMA(66), Z => n223);
   U66 : INVX0 port map( INP => RAMA(71), ZN => n18);
   U67 : INVX0 port map( INP => n18, ZN => n19);
   U68 : XOR2X1 port map( IN1 => n86, IN2 => RAMB(103), Q => addout_103_port);
   U69 : XOR2X1 port map( IN1 => RAMB(35), IN2 => n99, Q => addout_35_port);
   U70 : XOR2X1 port map( IN1 => RAMB(3), IN2 => n59, Q => addout_3_port);
   U71 : XOR2X1 port map( IN1 => RAMB(32), IN2 => n83, Q => addout_32_port);
   U72 : XOR2X1 port map( IN1 => RAMB(0), IN2 => n84, Q => addout_0_port);
   U73 : NBUFFX2 port map( INP => RAMA(127), Z => n28);
   U74 : XOR2X1 port map( IN1 => RAMB(49), IN2 => n51, Q => addout_49_port);
   U75 : XOR2X1 port map( IN1 => RAMB(54), IN2 => n54, Q => addout_54_port);
   U76 : XOR2X1 port map( IN1 => RAMB(1), IN2 => n130, Q => addout_1_port);
   U77 : NBUFFX2 port map( INP => RAMA(20), Z => n132);
   U78 : NBUFFX2 port map( INP => RAMA(113), Z => n57);
   U79 : NBUFFX2 port map( INP => RAMA(36), Z => n129);
   U80 : NBUFFX2 port map( INP => RAMA(69), Z => n109);
   U81 : NBUFFX2 port map( INP => RAMA(5), Z => n60);
   U82 : NBUFFX2 port map( INP => RAMA(47), Z => n134);
   U83 : NBUFFX2 port map( INP => RAMA(90), Z => n123);
   U84 : NBUFFX2 port map( INP => RAMA(65), Z => n49);
   U85 : NBUFFX2 port map( INP => RAMA(27), Z => n68);
   U86 : NBUFFX2 port map( INP => RAMA(87), Z => n77);
   U87 : NBUFFX2 port map( INP => RAMA(12), Z => n75);
   U88 : NBUFFX2 port map( INP => RAMA(50), Z => n116);
   U89 : NBUFFX2 port map( INP => RAMA(11), Z => n97);
   U90 : INVX0 port map( INP => n20, ZN => n21);
   U91 : NBUFFX2 port map( INP => RAMA(18), Z => n55);
   U92 : NBUFFX2 port map( INP => RAMA(7), Z => n111);
   U93 : NBUFFX2 port map( INP => RAMA(96), Z => n114);
   U94 : INVX0 port map( INP => RAMA(84), ZN => n32);
   U95 : XOR2X1 port map( IN1 => n1177, IN2 => n140, Q => addout_33_port);
   U96 : NBUFFX2 port map( INP => RAMA(23), Z => n43);
   U97 : NBUFFX2 port map( INP => RAMA(39), Z => n64);
   U98 : NBUFFX2 port map( INP => RAMA(107), Z => n87);
   U99 : NBUFFX2 port map( INP => RAMA(55), Z => n69);
   U100 : NBUFFX2 port map( INP => RAMA(79), Z => n115);
   U101 : NBUFFX2 port map( INP => RAMA(58), Z => n124);
   U102 : NBUFFX2 port map( INP => RAMA(60), Z => n81);
   U103 : NBUFFX2 port map( INP => RAMA(31), Z => n98);
   U104 : NBUFFX2 port map( INP => RAMA(101), Z => n94);
   U105 : NBUFFX2 port map( INP => RAMA(83), Z => n63);
   U106 : NBUFFX2 port map( INP => RAMA(6), Z => n135);
   U107 : NBUFFX2 port map( INP => RAMA(114), Z => n103);
   U108 : NBUFFX2 port map( INP => RAMA(118), Z => n80);
   U109 : INVX0 port map( INP => RAMA(85), ZN => n90);
   U110 : NBUFFX2 port map( INP => RAMA(119), Z => n47);
   U111 : NBUFFX2 port map( INP => RAMA(34), Z => n108);
   U112 : NBUFFX2 port map( INP => RAMA(86), Z => n95);
   U113 : NBUFFX2 port map( INP => RAMA(63), Z => n78);
   U114 : INVX0 port map( INP => RAMA(100), ZN => n142);
   U115 : NBUFFX2 port map( INP => RAMA(4), Z => n89);
   U116 : NBUFFX2 port map( INP => RAMA(75), Z => n42);
   U117 : NBUFFX2 port map( INP => RAMA(38), Z => n120);
   U118 : NBUFFX2 port map( INP => RAMA(35), Z => n99);
   U119 : NBUFFX2 port map( INP => RAMA(78), Z => n107);
   U120 : NBUFFX2 port map( INP => RAMA(46), Z => n85);
   U121 : INVX0 port map( INP => RAMA(98), ZN => n22);
   U122 : INVX0 port map( INP => n22, ZN => n23);
   U123 : INVX0 port map( INP => RAMA(116), ZN => n29);
   U124 : NBUFFX2 port map( INP => RAMA(111), Z => n41);
   U125 : NBUFFX2 port map( INP => RAMA(3), Z => n59);
   U126 : NBUFFX2 port map( INP => RAMA(103), Z => n86);
   U127 : AND2X4 port map( IN1 => RAMB(104), IN2 => RAMA(104), Q => 
                           andout_104_port);
   U128 : NBUFFX2 port map( INP => RAMA(14), Z => n125);
   U129 : NBUFFX2 port map( INP => RAMA(32), Z => n83);
   U130 : NBUFFX2 port map( INP => RAMA(49), Z => n51);
   U131 : NBUFFX2 port map( INP => RAMA(67), Z => n79);
   U132 : NBUFFX2 port map( INP => RAMA(54), Z => n54);
   U133 : NBUFFX2 port map( INP => RAMA(64), Z => n121);
   U134 : NBUFFX2 port map( INP => RAMA(51), Z => n133);
   U135 : NBUFFX2 port map( INP => RAMA(1), Z => n130);
   U136 : NBUFFX2 port map( INP => RAMA(15), Z => n101);
   U137 : NBUFFX2 port map( INP => RAMA(81), Z => n118);
   U138 : NBUFFX2 port map( INP => RAMA(17), Z => n122);
   U139 : NBUFFX2 port map( INP => RAMA(29), Z => n126);
   U140 : NBUFFX2 port map( INP => RAMA(62), Z => n52);
   U141 : NBUFFX2 port map( INP => RAMA(59), Z => n53);
   U142 : NBUFFX2 port map( INP => RAMA(76), Z => n137);
   U143 : NBUFFX2 port map( INP => RAMA(102), Z => n88);
   U144 : NBUFFX2 port map( INP => RAMA(0), Z => n84);
   U145 : NBUFFX2 port map( INP => RAMA(9), Z => n92);
   U146 : INVX0 port map( INP => RAMA(91), ZN => n70);
   U147 : NBUFFX2 port map( INP => RAMA(28), Z => n119);
   U148 : INVX0 port map( INP => RAMA(97), ZN => n24);
   U149 : INVX0 port map( INP => n24, ZN => n25);
   U150 : NBUFFX2 port map( INP => RAMA(70), Z => n58);
   U151 : NBUFFX2 port map( INP => RAMA(53), Z => n131);
   U152 : NBUFFX2 port map( INP => RAMA(19), Z => n72);
   U153 : NBUFFX2 port map( INP => RAMA(82), Z => n105);
   U154 : NBUFFX2 port map( INP => RAMA(77), Z => n62);
   U155 : INVX0 port map( INP => RAMA(117), ZN => n45);
   U156 : IBUFFX16 port map( INP => RAMA(95), ZN => n211);
   U157 : INVX0 port map( INP => RAMA(104), ZN => n202);
   U158 : XNOR2X2 port map( IN1 => RAMA(105), IN2 => n1249, Q => 
                           addout_105_port);
   U159 : INVX0 port map( INP => RAMA(126), ZN => n214);
   U160 : AO22X1 port map( IN1 => n995, IN2 => andout_48_port, IN3 => n996, IN4
                           => addout_48_port, Q => n703);
   U161 : INVX0 port map( INP => RAMA(74), ZN => n138);
   U162 : NBUFFX2 port map( INP => RAMA(115), Z => n26);
   U163 : XNOR2X2 port map( IN1 => RAMA(110), IN2 => n1254, Q => 
                           addout_110_port);
   U164 : XOR2X1 port map( IN1 => RAMB(48), IN2 => n1, Q => addout_48_port);
   U165 : INVX0 port map( INP => RAMA(33), ZN => n140);
   U166 : INVX0 port map( INP => n138, ZN => n27);
   U167 : INVX0 port map( INP => n29, ZN => n30);
   U168 : INVX0 port map( INP => n32, ZN => n33);
   U169 : XOR2X1 port map( IN1 => RAMB(116), IN2 => n30, Q => addout_116_port);
   U170 : INVX0 port map( INP => n200, ZN => n35);
   U171 : AND2X4 port map( IN1 => RAMB(24), IN2 => n36, Q => andout_24_port);
   U172 : IBUFFX16 port map( INP => RAMA(93), ZN => n38);
   U173 : INVX0 port map( INP => n38, ZN => n39);
   U174 : XOR2X1 port map( IN1 => RAMB(84), IN2 => n33, Q => addout_84_port);
   U175 : DELLN1X2 port map( INP => RAMA(44), Z => n44);
   U176 : INVX0 port map( INP => n45, ZN => n46);
   U177 : AND2X4 port map( IN1 => RAMB(119), IN2 => n47, Q => andout_119_port);
   U311 : AND2X4 port map( IN1 => RAMB(65), IN2 => n49, Q => andout_65_port);
   U312 : AND2X4 port map( IN1 => RAMB(59), IN2 => n53, Q => andout_59_port);
   U313 : AND2X4 port map( IN1 => RAMB(80), IN2 => n56, Q => andout_80_port);
   U314 : AND2X4 port map( IN1 => RAMB(113), IN2 => n57, Q => andout_113_port);
   U315 : DELLN1X2 port map( INP => RAMA(41), Z => n61);
   U317 : INVX0 port map( INP => n65, ZN => n66);
   U318 : AND2X4 port map( IN1 => RAMB(5), IN2 => n60, Q => andout_5_port);
   U320 : AND2X4 port map( IN1 => RAMB(3), IN2 => n59, Q => andout_3_port);
   U321 : INVX0 port map( INP => n70, ZN => n71);
   U322 : AND2X4 port map( IN1 => RAMB(27), IN2 => n68, Q => andout_27_port);
   U323 : AND2X4 port map( IN1 => RAMB(55), IN2 => n69, Q => andout_55_port);
   U325 : AND2X4 port map( IN1 => RAMB(25), IN2 => n73, Q => andout_25_port);
   U326 : DELLN1X2 port map( INP => RAMA(125), Z => n76);
   U327 : AND2X4 port map( IN1 => RAMB(125), IN2 => n76, Q => andout_125_port);
   U328 : AND2X4 port map( IN1 => RAMB(87), IN2 => n77, Q => andout_87_port);
   U329 : AND2X4 port map( IN1 => RAMB(52), IN2 => n31, Q => andout_52_port);
   U330 : AND2X4 port map( IN1 => RAMB(48), IN2 => n21, Q => andout_48_port);
   U331 : AND2X4 port map( IN1 => RAMB(63), IN2 => n78, Q => andout_63_port);
   U332 : AND2X4 port map( IN1 => RAMB(40), IN2 => n74, Q => andout_40_port);
   U333 : AND2X4 port map( IN1 => RAMB(12), IN2 => n75, Q => andout_12_port);
   U334 : AND2X4 port map( IN1 => RAMB(67), IN2 => n79, Q => andout_67_port);
   U335 : AND2X4 port map( IN1 => RAMB(118), IN2 => n80, Q => andout_118_port);
   U336 : AND2X4 port map( IN1 => RAMB(46), IN2 => n85, Q => andout_46_port);
   U337 : AND2X4 port map( IN1 => RAMB(42), IN2 => n82, Q => andout_42_port);
   U338 : AND2X4 port map( IN1 => RAMB(32), IN2 => n83, Q => andout_32_port);
   U340 : AND2X4 port map( IN1 => RAMB(0), IN2 => n84, Q => andout_0_port);
   U341 : AND2X4 port map( IN1 => RAMB(107), IN2 => n87, Q => andout_107_port);
   U342 : AND2X4 port map( IN1 => RAMB(102), IN2 => n88, Q => andout_102_port);
   U343 : INVX0 port map( INP => n90, ZN => n91);
   U344 : AND2X4 port map( IN1 => RAMB(98), IN2 => n23, Q => andout_98_port);
   U345 : AND2X4 port map( IN1 => RAMB(11), IN2 => n97, Q => andout_11_port);
   U346 : AND2X4 port map( IN1 => RAMB(61), IN2 => n100, Q => andout_61_port);
   U347 : AND2X4 port map( IN1 => RAMB(114), IN2 => n103, Q => andout_114_port)
                           ;
   U349 : AND2X4 port map( IN1 => RAMB(8), IN2 => n102, Q => andout_8_port);
   U350 : AND2X4 port map( IN1 => RAMB(15), IN2 => n101, Q => andout_15_port);
   U351 : AND2X4 port map( IN1 => RAMB(106), IN2 => n106, Q => andout_106_port)
                           ;
   U352 : AND2X4 port map( IN1 => RAMB(78), IN2 => n107, Q => andout_78_port);
   U353 : AND2X4 port map( IN1 => RAMB(69), IN2 => n109, Q => andout_69_port);
   U354 : AND2X4 port map( IN1 => RAMB(7), IN2 => n111, Q => andout_7_port);
   U355 : INVX0 port map( INP => n112, ZN => n113);
   U356 : AND2X4 port map( IN1 => RAMB(37), IN2 => n48, Q => andout_37_port);
   U357 : AND2X4 port map( IN1 => RAMB(50), IN2 => n116, Q => andout_50_port);
   U358 : AND2X4 port map( IN1 => RAMB(35), IN2 => n99, Q => andout_35_port);
   U359 : AND2X4 port map( IN1 => RAMB(64), IN2 => n121, Q => andout_64_port);
   U360 : AND2X4 port map( IN1 => RAMB(17), IN2 => n122, Q => andout_17_port);
   U361 : AND2X4 port map( IN1 => RAMB(120), IN2 => n2, Q => andout_120_port);
   U362 : AND2X4 port map( IN1 => RAMB(13), IN2 => n127, Q => andout_13_port);
   U363 : AND2X4 port map( IN1 => n17, IN2 => n129, Q => andout_36_port);
   U364 : AND2X4 port map( IN1 => RAMB(1), IN2 => n130, Q => andout_1_port);
   U365 : AND2X4 port map( IN1 => RAMB(41), IN2 => n61, Q => andout_41_port);
   U366 : AND2X4 port map( IN1 => RAMB(116), IN2 => n30, Q => andout_116_port);
   U367 : AND2X4 port map( IN1 => RAMB(20), IN2 => n132, Q => andout_20_port);
   U368 : AND2X4 port map( IN1 => RAMB(43), IN2 => n40, Q => andout_43_port);
   U369 : AND2X4 port map( IN1 => RAMB(51), IN2 => n133, Q => andout_51_port);
   U370 : AND2X4 port map( IN1 => RAMB(56), IN2 => n136, Q => andout_56_port);
   U371 : AND2X4 port map( IN1 => RAMB(6), IN2 => n135, Q => andout_6_port);
   U372 : AND2X4 port map( IN1 => RAMB(99), IN2 => n34, Q => andout_99_port);
   U373 : XOR2X1 port map( IN1 => RAMB(23), IN2 => n43, Q => addout_23_port);
   U374 : AND2X4 port map( IN1 => RAMB(23), IN2 => n43, Q => andout_23_port);
   U375 : AND2X4 port map( IN1 => RAMB(62), IN2 => n52, Q => andout_62_port);
   U376 : AND2X4 port map( IN1 => RAMB(76), IN2 => n137, Q => andout_76_port);
   U377 : AND2X4 port map( IN1 => RAMB(19), IN2 => n72, Q => andout_19_port);
   U378 : AND2X4 port map( IN1 => RAMB(111), IN2 => n41, Q => andout_111_port);
   U379 : AND2X4 port map( IN1 => RAMB(83), IN2 => n63, Q => andout_83_port);
   U380 : AND2X4 port map( IN1 => RAMB(86), IN2 => n95, Q => andout_86_port);
   U381 : AND2X4 port map( IN1 => RAMB(31), IN2 => n98, Q => andout_31_port);
   U382 : XNOR2X2 port map( IN1 => n23, IN2 => n161, Q => add_rnd_const_98_port
                           );
   U383 : AND2X4 port map( IN1 => RAMB(77), IN2 => n62, Q => andout_77_port);
   U385 : AND2X4 port map( IN1 => RAMB(60), IN2 => n81, Q => andout_60_port);
   U386 : AND2X4 port map( IN1 => RAMB(9), IN2 => n92, Q => andout_9_port);
   U387 : AND2X4 port map( IN1 => RAMB(10), IN2 => n93, Q => andout_10_port);
   U389 : XNOR2X2 port map( IN1 => n4, IN2 => n163, Q => add_rnd_const_105_port
                           );
   U390 : AND2X4 port map( IN1 => RAMB(105), IN2 => n4, Q => andout_105_port);
   U391 : AND2X4 port map( IN1 => RAMB(73), IN2 => n110, Q => andout_73_port);
   U393 : AND2X4 port map( IN1 => RAMB(54), IN2 => n54, Q => andout_54_port);
   U394 : AND2X4 port map( IN1 => RAMB(72), IN2 => n128, Q => andout_72_port);
   U395 : AND2X4 port map( IN1 => RAMB(16), IN2 => n117, Q => andout_16_port);
   U398 : AND2X4 port map( IN1 => RAMB(28), IN2 => n119, Q => andout_28_port);
   U399 : AND2X4 port map( IN1 => RAMB(47), IN2 => n134, Q => andout_47_port);
   U400 : AND2X4 port map( IN1 => RAMB(82), IN2 => n105, Q => andout_82_port);
   U401 : INVX0 port map( INP => n138, ZN => n139);
   U402 : INVX0 port map( INP => n140, ZN => n141);
   U403 : AND2X4 port map( IN1 => RAMB(97), IN2 => n25, Q => andout_97_port);
   U404 : AND2X4 port map( IN1 => RAMB(117), IN2 => n46, Q => andout_117_port);
   U405 : XOR2X1 port map( IN1 => RAMB(44), IN2 => n44, Q => addout_44_port);
   U406 : NAND2X0 port map( IN1 => n953, IN2 => n9, QN => perm_output(7));
   U407 : AND2X4 port map( IN1 => RAMB(30), IN2 => n37, Q => andout_30_port);
   U408 : AND2X4 port map( IN1 => n16, IN2 => n64, Q => andout_39_port);
   U409 : AND2X4 port map( IN1 => RAMB(44), IN2 => n44, Q => andout_44_port);
   U410 : AND2X4 port map( IN1 => RAMB(34), IN2 => n108, Q => andout_34_port);
   U411 : AND2X4 port map( IN1 => RAMB(14), IN2 => n125, Q => andout_14_port);
   U413 : AND2X4 port map( IN1 => RAMB(29), IN2 => n126, Q => andout_29_port);
   U414 : INVX0 port map( INP => n142, ZN => n143);
   U415 : AND2X4 port map( IN1 => RAMB(100), IN2 => n143, Q => andout_100_port)
                           ;
   U416 : AND2X4 port map( IN1 => RAMB(38), IN2 => n120, Q => andout_38_port);
   U417 : AND2X4 port map( IN1 => RAMB(45), IN2 => n67, Q => andout_45_port);
   U418 : AND2X4 port map( IN1 => RAMB(71), IN2 => n19, Q => andout_71_port);
   U419 : AND2X4 port map( IN1 => RAMB(4), IN2 => n89, Q => andout_4_port);
   U420 : AND2X4 port map( IN1 => RAMB(96), IN2 => n114, Q => andout_96_port);
   U422 : AND2X4 port map( IN1 => RAMB(110), IN2 => RAMA(110), Q => 
                           andout_110_port);
   U423 : AND2X4 port map( IN1 => RAMB(49), IN2 => n51, Q => andout_49_port);
   U424 : XOR2X1 port map( IN1 => n1239, IN2 => n211, Q => addout_95_port);
   U425 : AND2X4 port map( IN1 => RAMB(18), IN2 => n55, Q => andout_18_port);
   U426 : AND2X4 port map( IN1 => RAMB(68), IN2 => n220, Q => andout_68_port);
   U427 : XOR2X1 port map( IN1 => RAMB(85), IN2 => n91, Q => addout_85_port);
   U428 : INVX0 port map( INP => n202, ZN => n144);
   U430 : AND2X4 port map( IN1 => RAMB(53), IN2 => n131, Q => andout_53_port);
   U431 : INVX0 port map( INP => n200, ZN => n201);
   U432 : INVX0 port map( INP => n202, ZN => n203);
   U433 : NAND2X0 port map( IN1 => n467, IN2 => n11, QN => perm_output(88));
   U434 : AND2X4 port map( IN1 => RAMB(112), IN2 => n8, Q => andout_112_port);
   U435 : AND2X4 port map( IN1 => RAMB(75), IN2 => n42, Q => andout_75_port);
   U436 : NBUFFX2 port map( INP => RAMA(26), Z => n205);
   U437 : AND2X4 port map( IN1 => RAMB(101), IN2 => n94, Q => andout_101_port);
   U438 : AND2X4 port map( IN1 => RAMB(91), IN2 => n71, Q => andout_91_port);
   U441 : AND2X4 port map( IN1 => RAMB(90), IN2 => n123, Q => andout_90_port);
   U442 : NAND2X0 port map( IN1 => n653, IN2 => n12, QN => perm_output(57));
   U444 : AND2X4 port map( IN1 => RAMB(89), IN2 => n66, Q => andout_89_port);
   U446 : NBUFFX2 port map( INP => RAMA(2), Z => n208);
   U447 : AND2X4 port map( IN1 => RAMB(124), IN2 => n50, Q => andout_124_port);
   U452 : AND2X4 port map( IN1 => RAMB(70), IN2 => n58, Q => andout_70_port);
   U455 : AND2X4 port map( IN1 => RAMB(84), IN2 => n33, Q => andout_84_port);
   U456 : INVX0 port map( INP => n209, ZN => n204);
   U470 : INVX0 port map( INP => RAMA(22), ZN => n209);
   U474 : NBUFFX2 port map( INP => RAMA(108), Z => n213);
   U476 : XOR2X1 port map( IN1 => RAMB(26), IN2 => n205, Q => addout_26_port);
   U483 : IBUFFX16 port map( INP => RAMA(57), ZN => n206);
   U486 : INVX0 port map( INP => n206, ZN => n207);
   U489 : INVX0 port map( INP => n209, ZN => n210);
   U495 : XOR2X1 port map( IN1 => RAMB(2), IN2 => n208, Q => addout_2_port);
   U496 : INVX0 port map( INP => n211, ZN => n212);
   U500 : XOR2X1 port map( IN1 => RAMB(22), IN2 => n204, Q => addout_22_port);
   U505 : XOR2X1 port map( IN1 => RAMB(108), IN2 => n213, Q => addout_108_port)
                           ;
   U506 : XOR2X1 port map( IN1 => n1232, IN2 => n216, Q => addout_88_port);
   U509 : NAND2X0 port map( IN1 => n863, IN2 => n15, QN => perm_output(22));
   U510 : NBUFFX2 port map( INP => RAMA(92), Z => n218);
   U512 : NBUFFX2 port map( INP => RAMA(121), Z => n219);
   U513 : XOR2X1 port map( IN1 => n1267, IN2 => n221, Q => addout_123_port);
   U516 : NBUFFX2 port map( INP => RAMA(68), Z => n220);
   U520 : AND2X4 port map( IN1 => RAMB(85), IN2 => n91, Q => andout_85_port);
   U523 : AND2X4 port map( IN1 => RAMB(81), IN2 => n118, Q => andout_81_port);
   U524 : INVX0 port map( INP => n214, ZN => n215);
   U527 : INVX0 port map( INP => n216, ZN => n217);
   U537 : XOR2X1 port map( IN1 => RAMB(126), IN2 => n215, Q => addout_126_port)
                           ;
   U540 : NAND2X0 port map( IN1 => n245, IN2 => n10, QN => perm_output(125));
   U542 : NBUFFX2 port map( INP => n1005, Z => n1129);
   U547 : XOR2X1 port map( IN1 => RAMB(121), IN2 => n219, Q => addout_121_port)
                           ;
   U548 : XOR2X1 port map( IN1 => RAMB(92), IN2 => n218, Q => addout_92_port);
   U552 : XOR2X1 port map( IN1 => RAMB(68), IN2 => n220, Q => addout_68_port);
   U554 : AND2X4 port map( IN1 => RAMB(57), IN2 => RAMA(57), Q => 
                           andout_57_port);
   U556 : AND2X4 port map( IN1 => RAMB(127), IN2 => n28, Q => andout_127_port);
   U557 : AND2X4 port map( IN1 => RAMB(122), IN2 => n96, Q => andout_122_port);
   U560 : IBUFFX16 port map( INP => RAMA(123), ZN => n221);
   U562 : INVX0 port map( INP => n221, ZN => n222);
   U565 : AND2X4 port map( IN1 => RAMB(94), IN2 => n113, Q => andout_94_port);
   U566 : XOR2X1 port map( IN1 => RAMB(93), IN2 => n39, Q => addout_93_port);
   U569 : NAND2X0 port map( IN1 => n233, IN2 => n14, QN => perm_output(127));
   U570 : NAND2X0 port map( IN1 => n545, IN2 => n13, QN => perm_output(75));
   U571 : AND2X4 port map( IN1 => RAMB(93), IN2 => n39, Q => andout_93_port);
   U608 : AND2X4 port map( IN1 => RAMB(79), IN2 => n115, Q => andout_79_port);
   U609 : AND2X4 port map( IN1 => RAMB(58), IN2 => n124, Q => andout_58_port);
   U610 : NAND2X0 port map( IN1 => n179, IN2 => n152, QN => n183);
   U611 : NAND2X0 port map( IN1 => n152, IN2 => n1143, QN => n188);
   U612 : NAND2X0 port map( IN1 => n1143, IN2 => instruction_10_port, QN => 
                           n145);
   U613 : NAND2X0 port map( IN1 => n187, IN2 => n1143, QN => n150);
   U614 : NAND2X0 port map( IN1 => n1274, IN2 => n1275, QN => n155);
   U615 : NBUFFX2 port map( INP => n1003, Z => n1111);
   U616 : NBUFFX2 port map( INP => n1003, Z => n1112);
   U617 : NBUFFX2 port map( INP => n1003, Z => n1113);
   U618 : NBUFFX2 port map( INP => n1003, Z => n1114);
   U619 : NBUFFX2 port map( INP => n1003, Z => n1115);
   U620 : NBUFFX2 port map( INP => n1003, Z => n1116);
   U621 : NBUFFX2 port map( INP => n1003, Z => n1117);
   U622 : NBUFFX2 port map( INP => n1003, Z => n1118);
   U623 : NBUFFX2 port map( INP => n1003, Z => n1119);
   U624 : NBUFFX2 port map( INP => n1003, Z => n1120);
   U625 : NBUFFX2 port map( INP => n994, Z => n1045);
   U626 : NBUFFX2 port map( INP => n994, Z => n1046);
   U627 : NBUFFX2 port map( INP => n994, Z => n1047);
   U628 : NBUFFX2 port map( INP => n994, Z => n1048);
   U629 : NBUFFX2 port map( INP => n994, Z => n1049);
   U630 : NBUFFX2 port map( INP => n994, Z => n1050);
   U631 : NBUFFX2 port map( INP => n994, Z => n1051);
   U632 : NBUFFX2 port map( INP => n994, Z => n1052);
   U633 : NBUFFX2 port map( INP => n994, Z => n1053);
   U634 : NBUFFX2 port map( INP => n994, Z => n1054);
   U635 : NBUFFX2 port map( INP => n990, Z => n1012);
   U636 : NBUFFX2 port map( INP => n990, Z => n1013);
   U637 : NBUFFX2 port map( INP => n990, Z => n1014);
   U638 : NBUFFX2 port map( INP => n990, Z => n1015);
   U639 : NBUFFX2 port map( INP => n990, Z => n1016);
   U640 : NBUFFX2 port map( INP => n990, Z => n1017);
   U641 : NBUFFX2 port map( INP => n990, Z => n1018);
   U642 : NBUFFX2 port map( INP => n990, Z => n1019);
   U643 : NBUFFX2 port map( INP => n990, Z => n1020);
   U644 : NBUFFX2 port map( INP => n990, Z => n1021);
   U645 : NBUFFX2 port map( INP => n991, Z => n1023);
   U646 : NBUFFX2 port map( INP => n991, Z => n1024);
   U647 : NBUFFX2 port map( INP => n991, Z => n1025);
   U648 : NBUFFX2 port map( INP => n991, Z => n1026);
   U649 : NBUFFX2 port map( INP => n991, Z => n1027);
   U650 : NBUFFX2 port map( INP => n991, Z => n1028);
   U651 : NBUFFX2 port map( INP => n991, Z => n1029);
   U652 : NBUFFX2 port map( INP => n991, Z => n1030);
   U653 : NBUFFX2 port map( INP => n991, Z => n1031);
   U654 : NBUFFX2 port map( INP => n991, Z => n1032);
   U655 : NBUFFX2 port map( INP => n996, Z => n1067);
   U656 : NBUFFX2 port map( INP => n996, Z => n1068);
   U657 : NBUFFX2 port map( INP => n996, Z => n1069);
   U658 : NBUFFX2 port map( INP => n996, Z => n1070);
   U659 : NBUFFX2 port map( INP => n996, Z => n1071);
   U660 : NBUFFX2 port map( INP => n996, Z => n1072);
   U661 : NBUFFX2 port map( INP => n996, Z => n1073);
   U662 : NBUFFX2 port map( INP => n996, Z => n1074);
   U663 : NBUFFX2 port map( INP => n996, Z => n1075);
   U664 : NBUFFX2 port map( INP => n996, Z => n1076);
   U665 : NBUFFX2 port map( INP => n1010, Z => n1140);
   U666 : NBUFFX2 port map( INP => n1010, Z => n1139);
   U667 : NBUFFX2 port map( INP => n1010, Z => n1138);
   U668 : NBUFFX2 port map( INP => n1010, Z => n1137);
   U669 : NBUFFX2 port map( INP => n1010, Z => n1136);
   U670 : NBUFFX2 port map( INP => n1010, Z => n1135);
   U671 : NBUFFX2 port map( INP => n1010, Z => n1134);
   U672 : NBUFFX2 port map( INP => n1010, Z => n1133);
   U673 : NBUFFX2 port map( INP => n1010, Z => n1132);
   U674 : NBUFFX2 port map( INP => n1010, Z => n1131);
   U675 : NBUFFX2 port map( INP => n994, Z => n1044);
   U676 : NBUFFX2 port map( INP => n990, Z => n1011);
   U677 : NBUFFX2 port map( INP => n1003, Z => n1110);
   U678 : NBUFFX2 port map( INP => n991, Z => n1022);
   U679 : NBUFFX2 port map( INP => n996, Z => n1066);
   U680 : NBUFFX2 port map( INP => n1010, Z => n1130);
   U681 : NBUFFX2 port map( INP => n1005, Z => n1121);
   U682 : NBUFFX2 port map( INP => n1005, Z => n1122);
   U683 : NBUFFX2 port map( INP => n1005, Z => n1123);
   U684 : NBUFFX2 port map( INP => n1005, Z => n1124);
   U685 : NBUFFX2 port map( INP => n1005, Z => n1125);
   U686 : NBUFFX2 port map( INP => n1005, Z => n1126);
   U687 : NBUFFX2 port map( INP => n1005, Z => n1127);
   U688 : NBUFFX2 port map( INP => n1005, Z => n1128);
   U689 : NOR2X0 port map( IN1 => n1273, IN2 => n188, QN => ADDRA(3));
   U690 : INVX0 port map( INP => n148, ZN => n1273);
   U691 : NAND2X0 port map( IN1 => n1273, IN2 => n155, QN => n153);
   U692 : INVX0 port map( INP => n1142, ZN => n1278);
   U693 : INVX0 port map( INP => n188, ZN => n1280);
   U694 : NOR2X0 port map( IN1 => n1009, IN2 => n231, QN => n996);
   U695 : AND2X1 port map( IN1 => n226, IN2 => n1009, Q => n991);
   U696 : AND2X1 port map( IN1 => n225, IN2 => n1009, Q => n990);
   U697 : AND2X1 port map( IN1 => n227, IN2 => n1009, Q => n994);
   U698 : INVX0 port map( INP => instruction_9_port, ZN => n1008);
   U699 : INVX0 port map( INP => instruction_11_port, ZN => n1010);
   U700 : NBUFFX2 port map( INP => n998, Z => n1078);
   U701 : NBUFFX2 port map( INP => n998, Z => n1079);
   U702 : NBUFFX2 port map( INP => n998, Z => n1080);
   U703 : NBUFFX2 port map( INP => n998, Z => n1081);
   U704 : NBUFFX2 port map( INP => n998, Z => n1082);
   U705 : NBUFFX2 port map( INP => n998, Z => n1083);
   U706 : NBUFFX2 port map( INP => n998, Z => n1084);
   U707 : NBUFFX2 port map( INP => n998, Z => n1085);
   U708 : NBUFFX2 port map( INP => n998, Z => n1086);
   U709 : NBUFFX2 port map( INP => n998, Z => n1087);
   U710 : NBUFFX2 port map( INP => n995, Z => n1056);
   U711 : NBUFFX2 port map( INP => n995, Z => n1057);
   U712 : NBUFFX2 port map( INP => n995, Z => n1058);
   U713 : NBUFFX2 port map( INP => n995, Z => n1059);
   U714 : NBUFFX2 port map( INP => n995, Z => n1060);
   U715 : NBUFFX2 port map( INP => n995, Z => n1061);
   U716 : NBUFFX2 port map( INP => n995, Z => n1062);
   U717 : NBUFFX2 port map( INP => n995, Z => n1063);
   U718 : NBUFFX2 port map( INP => n995, Z => n1064);
   U719 : NBUFFX2 port map( INP => n995, Z => n1065);
   U720 : NBUFFX2 port map( INP => n999, Z => n1089);
   U721 : NBUFFX2 port map( INP => n999, Z => n1090);
   U722 : NBUFFX2 port map( INP => n999, Z => n1091);
   U723 : NBUFFX2 port map( INP => n999, Z => n1092);
   U724 : NBUFFX2 port map( INP => n999, Z => n1093);
   U725 : NBUFFX2 port map( INP => n999, Z => n1094);
   U726 : NBUFFX2 port map( INP => n999, Z => n1095);
   U727 : NBUFFX2 port map( INP => n999, Z => n1096);
   U728 : NBUFFX2 port map( INP => n999, Z => n1097);
   U729 : NBUFFX2 port map( INP => n999, Z => n1098);
   U730 : NBUFFX2 port map( INP => n1002, Z => n1100);
   U731 : NBUFFX2 port map( INP => n1002, Z => n1101);
   U732 : NBUFFX2 port map( INP => n1002, Z => n1102);
   U733 : NBUFFX2 port map( INP => n1002, Z => n1103);
   U734 : NBUFFX2 port map( INP => n1002, Z => n1104);
   U735 : NBUFFX2 port map( INP => n1002, Z => n1105);
   U736 : NBUFFX2 port map( INP => n1002, Z => n1106);
   U737 : NBUFFX2 port map( INP => n1002, Z => n1107);
   U738 : NBUFFX2 port map( INP => n1002, Z => n1108);
   U739 : NBUFFX2 port map( INP => n1002, Z => n1109);
   U740 : NBUFFX2 port map( INP => n993, Z => n1034);
   U741 : NBUFFX2 port map( INP => n993, Z => n1035);
   U742 : NBUFFX2 port map( INP => n993, Z => n1036);
   U743 : NBUFFX2 port map( INP => n993, Z => n1037);
   U744 : NBUFFX2 port map( INP => n993, Z => n1038);
   U745 : NBUFFX2 port map( INP => n993, Z => n1039);
   U746 : NBUFFX2 port map( INP => n993, Z => n1040);
   U747 : NBUFFX2 port map( INP => n993, Z => n1041);
   U748 : NBUFFX2 port map( INP => n993, Z => n1042);
   U749 : NBUFFX2 port map( INP => n993, Z => n1043);
   U750 : NBUFFX2 port map( INP => n998, Z => n1077);
   U751 : NBUFFX2 port map( INP => n995, Z => n1055);
   U752 : NBUFFX2 port map( INP => n999, Z => n1088);
   U753 : NBUFFX2 port map( INP => n1002, Z => n1099);
   U754 : NBUFFX2 port map( INP => n993, Z => n1033);
   U755 : INVX0 port map( INP => n155, ZN => n1272);
   U756 : NAND2X1 port map( IN1 => n160, IN2 => n1284, QN => n172);
   U757 : INVX0 port map( INP => n177, ZN => n1283);
   U758 : AND2X1 port map( IN1 => RAMB(121), IN2 => n219, Q => andout_121_port)
                           ;
   U759 : NOR2X0 port map( IN1 => n1274, IN2 => n1275, QN => n148);
   U760 : INVX0 port map( INP => RAMB(86), ZN => n1230);
   U761 : INVX0 port map( INP => RAMB(85), ZN => n1229);
   U762 : INVX0 port map( INP => RAMB(83), ZN => n1227);
   U763 : INVX0 port map( INP => RAMB(84), ZN => n1228);
   U764 : INVX0 port map( INP => RAMB(66), ZN => n1210);
   U765 : INVX0 port map( INP => RAMB(67), ZN => n1211);
   U766 : INVX0 port map( INP => RAMB(36), ZN => n1180);
   U767 : INVX0 port map( INP => RAMB(107), ZN => n1251);
   U768 : INVX0 port map( INP => RAMB(34), ZN => n1178);
   U769 : INVX0 port map( INP => RAMB(65), ZN => n1209);
   U770 : INVX0 port map( INP => RAMB(68), ZN => n1212);
   U771 : INVX0 port map( INP => RAMB(18), ZN => n1162);
   U772 : INVX0 port map( INP => RAMB(64), ZN => n1208);
   U773 : INVX0 port map( INP => RAMB(16), ZN => n1160);
   U774 : INVX0 port map( INP => RAMB(39), ZN => n1183);
   U775 : INVX0 port map( INP => RAMB(37), ZN => n1181);
   U776 : INVX0 port map( INP => RAMB(40), ZN => n1184);
   U777 : INVX0 port map( INP => RAMB(38), ZN => n1182);
   U778 : INVX0 port map( INP => RAMB(15), ZN => n1159);
   U779 : INVX0 port map( INP => RAMB(10), ZN => n1154);
   U780 : INVX0 port map( INP => RAMB(105), ZN => n1249);
   U781 : INVX0 port map( INP => RAMB(11), ZN => n1155);
   U782 : INVX0 port map( INP => RAMB(106), ZN => n1250);
   U783 : INVX0 port map( INP => RAMB(70), ZN => n1214);
   U784 : INVX0 port map( INP => RAMB(108), ZN => n1252);
   U785 : INVX0 port map( INP => RAMB(32), ZN => n1176);
   U786 : INVX0 port map( INP => RAMB(72), ZN => n1216);
   U787 : INVX0 port map( INP => RAMB(13), ZN => n1157);
   U788 : INVX0 port map( INP => RAMB(33), ZN => n1177);
   U789 : INVX0 port map( INP => RAMB(104), ZN => n1248);
   U790 : INVX0 port map( INP => RAMB(17), ZN => n1161);
   U791 : INVX0 port map( INP => RAMB(0), ZN => n1144);
   U792 : INVX0 port map( INP => RAMB(71), ZN => n1215);
   U793 : INVX0 port map( INP => RAMB(14), ZN => n1158);
   U794 : INVX0 port map( INP => RAMB(103), ZN => n1247);
   U795 : INVX0 port map( INP => RAMB(12), ZN => n1156);
   U796 : INVX0 port map( INP => RAMB(69), ZN => n1213);
   U797 : INVX0 port map( INP => RAMB(35), ZN => n1179);
   U798 : INVX0 port map( INP => RAMB(101), ZN => n1245);
   U799 : INVX0 port map( INP => RAMB(100), ZN => n1244);
   U800 : INVX0 port map( INP => RAMB(102), ZN => n1246);
   U801 : NAND2X0 port map( IN1 => n187, IN2 => n1278, QN => n194);
   U802 : INVX0 port map( INP => n146, ZN => n1277);
   U803 : INVX0 port map( INP => n150, ZN => n1279);
   U804 : INVX0 port map( INP => RAMB(58), ZN => n1202);
   U805 : INVX0 port map( INP => RAMB(97), ZN => n1241);
   U806 : INVX0 port map( INP => RAMB(98), ZN => n1242);
   U807 : INVX0 port map( INP => RAMB(90), ZN => n1234);
   U808 : INVX0 port map( INP => RAMB(87), ZN => n1231);
   U809 : INVX0 port map( INP => RAMB(94), ZN => n1238);
   U810 : INVX0 port map( INP => RAMB(9), ZN => n1153);
   U811 : INVX0 port map( INP => RAMB(55), ZN => n1199);
   U812 : INVX0 port map( INP => RAMB(23), ZN => n1167);
   U813 : INVX0 port map( INP => RAMB(24), ZN => n1168);
   U814 : INVX0 port map( INP => RAMB(93), ZN => n1237);
   U815 : INVX0 port map( INP => RAMB(91), ZN => n1235);
   U816 : INVX0 port map( INP => RAMB(88), ZN => n1232);
   U817 : INVX0 port map( INP => RAMB(56), ZN => n1200);
   U818 : INVX0 port map( INP => RAMB(57), ZN => n1201);
   U819 : INVX0 port map( INP => RAMB(59), ZN => n1203);
   U820 : INVX0 port map( INP => RAMB(96), ZN => n1240);
   U821 : INVX0 port map( INP => RAMB(62), ZN => n1206);
   U822 : INVX0 port map( INP => RAMB(6), ZN => n1150);
   U823 : INVX0 port map( INP => RAMB(95), ZN => n1239);
   U824 : INVX0 port map( INP => RAMB(7), ZN => n1151);
   U825 : INVX0 port map( INP => RAMB(2), ZN => n1146);
   U826 : INVX0 port map( INP => RAMB(126), ZN => n1270);
   U827 : INVX0 port map( INP => RAMB(8), ZN => n1152);
   U828 : INVX0 port map( INP => RAMB(61), ZN => n1205);
   U829 : INVX0 port map( INP => RAMB(125), ZN => n1269);
   U830 : INVX0 port map( INP => RAMB(123), ZN => n1267);
   U831 : INVX0 port map( INP => RAMB(127), ZN => n1271);
   U832 : INVX0 port map( INP => RAMB(92), ZN => n1236);
   U833 : INVX0 port map( INP => RAMB(63), ZN => n1207);
   U834 : INVX0 port map( INP => RAMB(60), ZN => n1204);
   U835 : INVX0 port map( INP => RAMB(124), ZN => n1268);
   U836 : INVX0 port map( INP => RAMB(5), ZN => n1149);
   U837 : INVX0 port map( INP => RAMB(89), ZN => n1233);
   U838 : INVX0 port map( INP => RAMB(4), ZN => n1148);
   U839 : INVX0 port map( INP => RAMB(3), ZN => n1147);
   U840 : INVX0 port map( INP => RAMB(99), ZN => n1243);
   U841 : INVX0 port map( INP => RAMB(29), ZN => n1173);
   U842 : INVX0 port map( INP => RAMB(76), ZN => n1220);
   U843 : INVX0 port map( INP => RAMB(19), ZN => n1163);
   U844 : INVX0 port map( INP => RAMB(26), ZN => n1170);
   U845 : INVX0 port map( INP => RAMB(28), ZN => n1172);
   U846 : INVX0 port map( INP => RAMB(30), ZN => n1174);
   U847 : INVX0 port map( INP => RAMB(21), ZN => n1165);
   U848 : INVX0 port map( INP => RAMB(50), ZN => n1194);
   U849 : INVX0 port map( INP => RAMB(27), ZN => n1171);
   U850 : INVX0 port map( INP => RAMB(80), ZN => n1224);
   U851 : INVX0 port map( INP => RAMB(49), ZN => n1193);
   U852 : INVX0 port map( INP => RAMB(51), ZN => n1195);
   U853 : INVX0 port map( INP => RAMB(25), ZN => n1169);
   U854 : INVX0 port map( INP => RAMB(20), ZN => n1164);
   U855 : INVX0 port map( INP => RAMB(48), ZN => n1192);
   U856 : INVX0 port map( INP => RAMB(78), ZN => n1222);
   U857 : INVX0 port map( INP => RAMB(1), ZN => n1145);
   U858 : INVX0 port map( INP => RAMB(81), ZN => n1225);
   U859 : INVX0 port map( INP => RAMB(53), ZN => n1197);
   U860 : INVX0 port map( INP => RAMB(82), ZN => n1226);
   U861 : INVX0 port map( INP => RAMB(22), ZN => n1166);
   U862 : INVX0 port map( INP => RAMB(45), ZN => n1189);
   U863 : INVX0 port map( INP => RAMB(54), ZN => n1198);
   U864 : INVX0 port map( INP => RAMB(119), ZN => n1263);
   U865 : INVX0 port map( INP => RAMB(42), ZN => n1186);
   U866 : INVX0 port map( INP => RAMB(47), ZN => n1191);
   U867 : INVX0 port map( INP => RAMB(41), ZN => n1185);
   U868 : INVX0 port map( INP => RAMB(77), ZN => n1221);
   U869 : INVX0 port map( INP => RAMB(79), ZN => n1223);
   U870 : INVX0 port map( INP => RAMB(43), ZN => n1187);
   U871 : INVX0 port map( INP => RAMB(114), ZN => n1258);
   U872 : INVX0 port map( INP => RAMB(73), ZN => n1217);
   U873 : INVX0 port map( INP => RAMB(46), ZN => n1190);
   U874 : INVX0 port map( INP => RAMB(74), ZN => n1218);
   U875 : INVX0 port map( INP => RAMB(75), ZN => n1219);
   U876 : INVX0 port map( INP => RAMB(31), ZN => n1175);
   U877 : INVX0 port map( INP => RAMB(112), ZN => n1256);
   U878 : INVX0 port map( INP => RAMB(113), ZN => n1257);
   U879 : INVX0 port map( INP => RAMB(52), ZN => n1196);
   U880 : INVX0 port map( INP => RAMB(110), ZN => n1254);
   U881 : INVX0 port map( INP => RAMB(111), ZN => n1255);
   U882 : INVX0 port map( INP => RAMB(109), ZN => n1253);
   U883 : INVX0 port map( INP => RAMB(122), ZN => n1266);
   U884 : INVX0 port map( INP => RAMB(44), ZN => n1188);
   U885 : INVX0 port map( INP => RAMB(115), ZN => n1259);
   U886 : INVX0 port map( INP => RAMB(121), ZN => n1265);
   U887 : INVX0 port map( INP => RAMB(116), ZN => n1260);
   U888 : INVX0 port map( INP => RAMB(118), ZN => n1262);
   U889 : INVX0 port map( INP => RAMB(117), ZN => n1261);
   U890 : INVX0 port map( INP => RAMB(120), ZN => n1264);
   U891 : INVX0 port map( INP => n1141, ZN => n1142);
   U892 : NOR2X0 port map( IN1 => n1277, IN2 => n152, QN => n193);
   U893 : INVX0 port map( INP => n186, ZN => n1276);
   U894 : NAND2X0 port map( IN1 => n1276, IN2 => n1281, QN => n192);
   U895 : INVX0 port map( INP => n1141, ZN => n1143);
   U896 : NOR2X0 port map( IN1 => n231, IN2 => instruction_8_port, QN => n993);
   U897 : NAND2X0 port map( IN1 => n148, IN2 => n1282, QN => n147);
   U898 : INVX0 port map( INP => instruction_8_port, ZN => n1009);
   U899 : AND2X1 port map( IN1 => n227, IN2 => instruction_8_port, Q => n995);
   U900 : AND2X1 port map( IN1 => n225, IN2 => instruction_8_port, Q => n999);
   U901 : AND2X1 port map( IN1 => n226, IN2 => instruction_8_port, Q => n998);
   U902 : NOR2X0 port map( IN1 => n1143, IN2 => n1273, QN => n154);
   U903 : INVX0 port map( INP => instruction_10_port, ZN => n1007);
   U904 : NAND2X1 port map( IN1 => n177, IN2 => n174, QN => n157);
   U905 : NOR2X0 port map( IN1 => n1287, IN2 => n1286, QN => n160);
   U906 : NAND2X0 port map( IN1 => ins_counter(0), IN2 => n199, QN => n197);
   U907 : NOR2X0 port map( IN1 => n1282, IN2 => ins_counter(3), QN => n152);
   U908 : NAND2X0 port map( IN1 => n194, IN2 => n188, QN => n196);
   U909 : NOR2X0 port map( IN1 => n1275, IN2 => ins_counter(0), QN => n179);
   U910 : INVX0 port map( INP => n160, ZN => n1285);
   U911 : NAND2X0 port map( IN1 => RNDCTR(2), IN2 => RNDCTR(0), QN => n161);
   U912 : NOR2X0 port map( IN1 => n1281, IN2 => ins_counter(4), QN => 
                           instruction_10_port);
   U913 : INVX0 port map( INP => ins_counter(1), ZN => n1275);
   U914 : INVX0 port map( INP => ins_counter(0), ZN => n1274);
   U915 : INVX0 port map( INP => ins_counter(4), ZN => n1282);
   U916 : NOR2X0 port map( IN1 => ins_counter(3), IN2 => ins_counter(4), QN => 
                           n187);
   U917 : NOR2X0 port map( IN1 => n1282, IN2 => ins_counter(1), QN => n186);
   U918 : NAND2X0 port map( IN1 => ins_counter(1), IN2 => instruction_10_port, 
                           QN => n146);
   U919 : NAND2X0 port map( IN1 => n160, IN2 => RNDCTR(0), QN => n159);
   U920 : INVX0 port map( INP => ins_counter(3), ZN => n1281);
   U921 : INVX0 port map( INP => ins_counter(2), ZN => n1141);
   U922 : INVX0 port map( INP => RNDCTR(0), ZN => n1284);
   U923 : NOR2X0 port map( IN1 => n1284, IN2 => RNDCTR(1), QN => n177);
   U924 : NOR2X0 port map( IN1 => RNDCTR(2), IN2 => RNDCTR(3), QN => n174);
   U925 : NAND2X1 port map( IN1 => RNDCTR(3), IN2 => n177, QN => n169);
   U926 : INVX0 port map( INP => RNDCTR(1), ZN => n1286);
   U927 : NAND2X1 port map( IN1 => RNDCTR(3), IN2 => n1284, QN => n164);
   U928 : INVX0 port map( INP => RNDCTR(2), ZN => n1287);
   U929 : NOR2X0 port map( IN1 => n1008, IN2 => n1007, QN => n227);
   U930 : NAND2X0 port map( IN1 => n1008, IN2 => n1007, QN => n231);
   U931 : NOR2X0 port map( IN1 => n1008, IN2 => instruction_10_port, QN => n226
                           );
   U932 : NOR2X0 port map( IN1 => n1007, IN2 => instruction_9_port, QN => n225)
                           ;
   U933 : AO22X1 port map( IN1 => eshift_127_port, IN2 => n1032, IN3 => n1021, 
                           IN4 => RAMB(116), Q => n224);
   U934 : AO221X1 port map( IN1 => n1271, IN2 => n1054, IN3 => n1043, IN4 => 
                           RAMB(127), IN5 => n224, Q => n230);
   U935 : AO22X1 port map( IN1 => addout_127_port, IN2 => n1076, IN3 => 
                           andout_127_port, IN4 => n1065, Q => n228);
   U936 : AO221X1 port map( IN1 => n28, IN2 => n1098, IN3 => n1087, IN4 => 
                           RAMB(31), IN5 => n228, Q => n229);
   U937 : OAI21X1 port map( IN1 => n230, IN2 => n229, IN3 => n1130, QN => n233)
                           ;
   U938 : OA22X1 port map( IN1 => n1270, IN2 => n1120, IN3 => n1199, IN4 => 
                           n1109, Q => n232);
   U939 : AO22X1 port map( IN1 => eshift_126_port, IN2 => n1032, IN3 => n1021, 
                           IN4 => RAMB(115), Q => n234);
   U940 : AO221X1 port map( IN1 => n1270, IN2 => n1054, IN3 => n1043, IN4 => 
                           RAMB(126), IN5 => n234, Q => n237);
   U941 : AO22X1 port map( IN1 => addout_126_port, IN2 => n1076, IN3 => 
                           andout_126_port, IN4 => n1065, Q => n235);
   U942 : AO221X1 port map( IN1 => n215, IN2 => n1098, IN3 => n1087, IN4 => 
                           RAMB(30), IN5 => n235, Q => n236);
   U943 : OAI21X1 port map( IN1 => n237, IN2 => n236, IN3 => n1130, QN => n239)
                           ;
   U944 : OA22X1 port map( IN1 => n1269, IN2 => n1120, IN3 => n1198, IN4 => 
                           n1109, Q => n238);
   U945 : NAND3X0 port map( IN1 => n239, IN2 => n1129, IN3 => n238, QN => 
                           perm_output(126));
   U946 : AO22X1 port map( IN1 => eshift_125_port, IN2 => n1032, IN3 => n1021, 
                           IN4 => RAMB(114), Q => n240);
   U947 : AO221X1 port map( IN1 => n1269, IN2 => n1054, IN3 => n1043, IN4 => 
                           RAMB(125), IN5 => n240, Q => n243);
   U948 : AO22X1 port map( IN1 => addout_125_port, IN2 => n1076, IN3 => 
                           andout_125_port, IN4 => n1065, Q => n241);
   U949 : AO221X1 port map( IN1 => n76, IN2 => n1098, IN3 => n1087, IN4 => 
                           RAMB(29), IN5 => n241, Q => n242);
   U950 : OAI21X1 port map( IN1 => n243, IN2 => n242, IN3 => n1130, QN => n245)
                           ;
   U951 : OA22X1 port map( IN1 => n1268, IN2 => n1120, IN3 => n1197, IN4 => 
                           n1109, Q => n244);
   U952 : AO22X1 port map( IN1 => eshift_124_port, IN2 => n1032, IN3 => n1021, 
                           IN4 => RAMB(113), Q => n246);
   U953 : AO221X1 port map( IN1 => n1268, IN2 => n1054, IN3 => n1043, IN4 => 
                           RAMB(124), IN5 => n246, Q => n249);
   U954 : AO22X1 port map( IN1 => addout_124_port, IN2 => n1076, IN3 => 
                           andout_124_port, IN4 => n1065, Q => n247);
   U955 : AO221X1 port map( IN1 => n50, IN2 => n1098, IN3 => n1087, IN4 => 
                           RAMB(28), IN5 => n247, Q => n248);
   U956 : OAI21X1 port map( IN1 => n249, IN2 => n248, IN3 => n1130, QN => n251)
                           ;
   U957 : OA22X1 port map( IN1 => n1267, IN2 => n1120, IN3 => n1196, IN4 => 
                           n1109, Q => n250);
   U958 : NAND3X0 port map( IN1 => n251, IN2 => n1129, IN3 => n250, QN => 
                           perm_output(124));
   U959 : AO22X1 port map( IN1 => eshift_123_port, IN2 => n1032, IN3 => n1021, 
                           IN4 => RAMB(112), Q => n252);
   U960 : AO221X1 port map( IN1 => n1267, IN2 => n1054, IN3 => n1043, IN4 => 
                           RAMB(123), IN5 => n252, Q => n255);
   U961 : AO22X1 port map( IN1 => addout_123_port, IN2 => n1076, IN3 => 
                           andout_123_port, IN4 => n1065, Q => n253);
   U962 : AO221X1 port map( IN1 => n222, IN2 => n1098, IN3 => n1087, IN4 => 
                           RAMB(27), IN5 => n253, Q => n254);
   U963 : OAI21X1 port map( IN1 => n255, IN2 => n254, IN3 => n1130, QN => n257)
                           ;
   U964 : OA22X1 port map( IN1 => n1266, IN2 => n1120, IN3 => n1195, IN4 => 
                           n1109, Q => n256);
   U965 : NAND3X0 port map( IN1 => n257, IN2 => n1129, IN3 => n256, QN => 
                           perm_output(123));
   U966 : AO22X1 port map( IN1 => eshift_122_port, IN2 => n1032, IN3 => n1021, 
                           IN4 => RAMB(111), Q => n258);
   U967 : AO221X1 port map( IN1 => n1266, IN2 => n1054, IN3 => n1043, IN4 => 
                           RAMB(122), IN5 => n258, Q => n261);
   U968 : AO22X1 port map( IN1 => addout_122_port, IN2 => n1076, IN3 => 
                           andout_122_port, IN4 => n1065, Q => n259);
   U969 : AO221X1 port map( IN1 => n96, IN2 => n1098, IN3 => n1087, IN4 => 
                           RAMB(26), IN5 => n259, Q => n260);
   U970 : OAI21X1 port map( IN1 => n261, IN2 => n260, IN3 => n1130, QN => n263)
                           ;
   U971 : OA22X1 port map( IN1 => n1265, IN2 => n1120, IN3 => n1194, IN4 => 
                           n1109, Q => n262);
   U972 : NAND3X0 port map( IN1 => n263, IN2 => n1129, IN3 => n262, QN => 
                           perm_output(122));
   U973 : AO22X1 port map( IN1 => eshift_121_port, IN2 => n1032, IN3 => n1021, 
                           IN4 => RAMB(110), Q => n264);
   U974 : AO221X1 port map( IN1 => n1265, IN2 => n1054, IN3 => n1043, IN4 => 
                           RAMB(121), IN5 => n264, Q => n267);
   U975 : AO22X1 port map( IN1 => addout_121_port, IN2 => n1076, IN3 => 
                           andout_121_port, IN4 => n1065, Q => n265);
   U976 : AO221X1 port map( IN1 => n219, IN2 => n1098, IN3 => n1087, IN4 => 
                           RAMB(25), IN5 => n265, Q => n266);
   U977 : OAI21X1 port map( IN1 => n267, IN2 => n266, IN3 => n1130, QN => n269)
                           ;
   U978 : OA22X1 port map( IN1 => n1264, IN2 => n1120, IN3 => n1193, IN4 => 
                           n1109, Q => n268);
   U979 : NAND3X0 port map( IN1 => n269, IN2 => n1129, IN3 => n268, QN => 
                           perm_output(121));
   U980 : AO22X1 port map( IN1 => eshift_120_port, IN2 => n1032, IN3 => n1021, 
                           IN4 => RAMB(109), Q => n270);
   U981 : AO221X1 port map( IN1 => n1264, IN2 => n1054, IN3 => n1043, IN4 => 
                           RAMB(120), IN5 => n270, Q => n273);
   U982 : AO22X1 port map( IN1 => addout_120_port, IN2 => n1076, IN3 => 
                           andout_120_port, IN4 => n1065, Q => n271);
   U983 : AO221X1 port map( IN1 => n2, IN2 => n1098, IN3 => n1087, IN4 => 
                           RAMB(24), IN5 => n271, Q => n272);
   U984 : OAI21X1 port map( IN1 => n273, IN2 => n272, IN3 => n1130, QN => n275)
                           ;
   U985 : OA22X1 port map( IN1 => n1263, IN2 => n1120, IN3 => n1192, IN4 => 
                           n1109, Q => n274);
   U986 : NAND3X0 port map( IN1 => n275, IN2 => n1129, IN3 => n274, QN => 
                           perm_output(120));
   U987 : AO22X1 port map( IN1 => eshift_119_port, IN2 => n1032, IN3 => n1021, 
                           IN4 => RAMB(108), Q => n276);
   U988 : AO221X1 port map( IN1 => n1263, IN2 => n1054, IN3 => n1043, IN4 => 
                           RAMB(119), IN5 => n276, Q => n279);
   U989 : AO22X1 port map( IN1 => addout_119_port, IN2 => n1076, IN3 => 
                           andout_119_port, IN4 => n1065, Q => n277);
   U990 : AO221X1 port map( IN1 => n47, IN2 => n1098, IN3 => n1087, IN4 => 
                           RAMB(23), IN5 => n277, Q => n278);
   U991 : OAI21X1 port map( IN1 => n279, IN2 => n278, IN3 => n1131, QN => n281)
                           ;
   U992 : OA22X1 port map( IN1 => n1262, IN2 => n1120, IN3 => n1191, IN4 => 
                           n1109, Q => n280);
   U993 : NAND3X0 port map( IN1 => n281, IN2 => n1129, IN3 => n280, QN => 
                           perm_output(119));
   U994 : AO22X1 port map( IN1 => eshift_118_port, IN2 => n1032, IN3 => n1021, 
                           IN4 => RAMB(107), Q => n282);
   U995 : AO221X1 port map( IN1 => n1262, IN2 => n1054, IN3 => n1043, IN4 => 
                           RAMB(118), IN5 => n282, Q => n285);
   U996 : AO22X1 port map( IN1 => addout_118_port, IN2 => n1076, IN3 => 
                           andout_118_port, IN4 => n1065, Q => n283);
   U997 : AO221X1 port map( IN1 => n80, IN2 => n1098, IN3 => n1087, IN4 => 
                           RAMB(22), IN5 => n283, Q => n284);
   U998 : OAI21X1 port map( IN1 => n285, IN2 => n284, IN3 => n1131, QN => n287)
                           ;
   U999 : OA22X1 port map( IN1 => n1261, IN2 => n1120, IN3 => n1190, IN4 => 
                           n1109, Q => n286);
   U1000 : NAND3X0 port map( IN1 => n287, IN2 => n1129, IN3 => n286, QN => 
                           perm_output(118));
   U1001 : AO22X1 port map( IN1 => eshift_117_port, IN2 => n1032, IN3 => n1021,
                           IN4 => RAMB(106), Q => n288);
   U1002 : AO221X1 port map( IN1 => n1261, IN2 => n1054, IN3 => n1043, IN4 => 
                           RAMB(117), IN5 => n288, Q => n291);
   U1003 : AO22X1 port map( IN1 => addout_117_port, IN2 => n1076, IN3 => 
                           andout_117_port, IN4 => n1065, Q => n289);
   U1004 : AO221X1 port map( IN1 => n46, IN2 => n1098, IN3 => n1087, IN4 => 
                           RAMB(21), IN5 => n289, Q => n290);
   U1005 : OAI21X1 port map( IN1 => n291, IN2 => n290, IN3 => n1131, QN => n293
                           );
   U1006 : OA22X1 port map( IN1 => n1260, IN2 => n1120, IN3 => n1189, IN4 => 
                           n1109, Q => n292);
   U1007 : NAND3X0 port map( IN1 => n293, IN2 => n1129, IN3 => n292, QN => 
                           perm_output(117));
   U1008 : AO22X1 port map( IN1 => eshift_116_port, IN2 => n1032, IN3 => n1021,
                           IN4 => RAMB(105), Q => n294);
   U1009 : AO221X1 port map( IN1 => n1260, IN2 => n1054, IN3 => n1043, IN4 => 
                           RAMB(116), IN5 => n294, Q => n297);
   U1010 : AO22X1 port map( IN1 => addout_116_port, IN2 => n1076, IN3 => 
                           andout_116_port, IN4 => n1065, Q => n295);
   U1011 : AO221X1 port map( IN1 => n30, IN2 => n1098, IN3 => n1087, IN4 => 
                           RAMB(20), IN5 => n295, Q => n296);
   U1012 : OAI21X1 port map( IN1 => n297, IN2 => n296, IN3 => n1131, QN => n299
                           );
   U1013 : OA22X1 port map( IN1 => n1259, IN2 => n1120, IN3 => n1188, IN4 => 
                           n1109, Q => n298);
   U1014 : NAND3X0 port map( IN1 => n299, IN2 => n1129, IN3 => n298, QN => 
                           perm_output(116));
   U1015 : AO22X1 port map( IN1 => eshift_115_port, IN2 => n1031, IN3 => n1020,
                           IN4 => RAMB(104), Q => n300);
   U1016 : AO221X1 port map( IN1 => n1259, IN2 => n1053, IN3 => n1042, IN4 => 
                           RAMB(115), IN5 => n300, Q => n303);
   U1017 : AO22X1 port map( IN1 => addout_115_port, IN2 => n1075, IN3 => 
                           andout_115_port, IN4 => n1064, Q => n301);
   U1018 : AO221X1 port map( IN1 => n26, IN2 => n1097, IN3 => n1086, IN4 => 
                           RAMB(19), IN5 => n301, Q => n302);
   U1019 : OAI21X1 port map( IN1 => n303, IN2 => n302, IN3 => n1131, QN => n305
                           );
   U1020 : OA22X1 port map( IN1 => n1258, IN2 => n1119, IN3 => n1187, IN4 => 
                           n1108, Q => n304);
   U1021 : NAND3X0 port map( IN1 => n305, IN2 => n1128, IN3 => n304, QN => 
                           perm_output(115));
   U1022 : AO22X1 port map( IN1 => eshift_114_port, IN2 => n1031, IN3 => n1020,
                           IN4 => RAMB(103), Q => n306);
   U1023 : AO221X1 port map( IN1 => n1258, IN2 => n1053, IN3 => n1042, IN4 => 
                           RAMB(114), IN5 => n306, Q => n309);
   U1024 : AO22X1 port map( IN1 => addout_114_port, IN2 => n1075, IN3 => 
                           andout_114_port, IN4 => n1064, Q => n307);
   U1025 : AO221X1 port map( IN1 => n103, IN2 => n1097, IN3 => n1086, IN4 => 
                           RAMB(18), IN5 => n307, Q => n308);
   U1026 : OAI21X1 port map( IN1 => n309, IN2 => n308, IN3 => n1131, QN => n311
                           );
   U1027 : OA22X1 port map( IN1 => n1257, IN2 => n1119, IN3 => n1186, IN4 => 
                           n1108, Q => n310);
   U1028 : NAND3X0 port map( IN1 => n311, IN2 => n1128, IN3 => n310, QN => 
                           perm_output(114));
   U1029 : AO22X1 port map( IN1 => eshift_113_port, IN2 => n1031, IN3 => n1020,
                           IN4 => RAMB(102), Q => n312);
   U1030 : AO221X1 port map( IN1 => n1257, IN2 => n1053, IN3 => n1042, IN4 => 
                           RAMB(113), IN5 => n312, Q => n315);
   U1031 : AO22X1 port map( IN1 => addout_113_port, IN2 => n1075, IN3 => 
                           andout_113_port, IN4 => n1064, Q => n313);
   U1032 : AO221X1 port map( IN1 => n57, IN2 => n1097, IN3 => n1086, IN4 => 
                           RAMB(17), IN5 => n313, Q => n314);
   U1033 : OAI21X1 port map( IN1 => n315, IN2 => n314, IN3 => n1131, QN => n317
                           );
   U1034 : OA22X1 port map( IN1 => n1256, IN2 => n1119, IN3 => n1185, IN4 => 
                           n1108, Q => n316);
   U1035 : NAND3X0 port map( IN1 => n317, IN2 => n1128, IN3 => n316, QN => 
                           perm_output(113));
   U1036 : AO22X1 port map( IN1 => eshift_112_port, IN2 => n1031, IN3 => n1020,
                           IN4 => RAMB(101), Q => n318);
   U1037 : AO221X1 port map( IN1 => n1256, IN2 => n1053, IN3 => n1042, IN4 => 
                           RAMB(112), IN5 => n318, Q => n321);
   U1038 : AO22X1 port map( IN1 => addout_112_port, IN2 => n1075, IN3 => 
                           andout_112_port, IN4 => n1064, Q => n319);
   U1039 : AO221X1 port map( IN1 => n8, IN2 => n1097, IN3 => n1086, IN4 => 
                           RAMB(16), IN5 => n319, Q => n320);
   U1040 : OAI21X1 port map( IN1 => n321, IN2 => n320, IN3 => n1131, QN => n323
                           );
   U1041 : OA22X1 port map( IN1 => n1255, IN2 => n1119, IN3 => n1184, IN4 => 
                           n1108, Q => n322);
   U1042 : NAND3X0 port map( IN1 => n323, IN2 => n1128, IN3 => n322, QN => 
                           perm_output(112));
   U1043 : AO22X1 port map( IN1 => eshift_111_port, IN2 => n1031, IN3 => n1020,
                           IN4 => RAMB(100), Q => n324);
   U1044 : AO221X1 port map( IN1 => n1255, IN2 => n1053, IN3 => n1042, IN4 => 
                           RAMB(111), IN5 => n324, Q => n327);
   U1045 : AO22X1 port map( IN1 => addout_111_port, IN2 => n1075, IN3 => 
                           andout_111_port, IN4 => n1064, Q => n325);
   U1046 : AO221X1 port map( IN1 => n41, IN2 => n1097, IN3 => n1086, IN4 => 
                           RAMB(15), IN5 => n325, Q => n326);
   U1047 : OAI21X1 port map( IN1 => n327, IN2 => n326, IN3 => n1131, QN => n329
                           );
   U1048 : OA22X1 port map( IN1 => n1254, IN2 => n1119, IN3 => n1183, IN4 => 
                           n1108, Q => n328);
   U1049 : NAND3X0 port map( IN1 => n329, IN2 => n1128, IN3 => n328, QN => 
                           perm_output(111));
   U1050 : AO22X1 port map( IN1 => eshift_110_port, IN2 => n1031, IN3 => n1020,
                           IN4 => RAMB(99), Q => n330);
   U1051 : AO221X1 port map( IN1 => n1254, IN2 => n1053, IN3 => n1042, IN4 => 
                           RAMB(110), IN5 => n330, Q => n333);
   U1052 : AO22X1 port map( IN1 => addout_110_port, IN2 => n1075, IN3 => 
                           andout_110_port, IN4 => n1064, Q => n331);
   U1053 : AO221X1 port map( IN1 => RAMA(110), IN2 => n1097, IN3 => n1086, IN4 
                           => RAMB(14), IN5 => n331, Q => n332);
   U1054 : OAI21X1 port map( IN1 => n333, IN2 => n332, IN3 => n1131, QN => n335
                           );
   U1055 : OA22X1 port map( IN1 => n1253, IN2 => n1119, IN3 => n1182, IN4 => 
                           n1108, Q => n334);
   U1056 : NAND3X0 port map( IN1 => n335, IN2 => n1128, IN3 => n334, QN => 
                           perm_output(110));
   U1057 : AO22X1 port map( IN1 => eshift_109_port, IN2 => n1031, IN3 => n1020,
                           IN4 => RAMB(98), Q => n336);
   U1058 : AO221X1 port map( IN1 => n1253, IN2 => n1053, IN3 => n1042, IN4 => 
                           RAMB(109), IN5 => n336, Q => n339);
   U1059 : AO22X1 port map( IN1 => addout_109_port, IN2 => n1075, IN3 => 
                           andout_109_port, IN4 => n1064, Q => n337);
   U1060 : AO221X1 port map( IN1 => n104, IN2 => n1097, IN3 => n1086, IN4 => 
                           RAMB(13), IN5 => n337, Q => n338);
   U1061 : OAI21X1 port map( IN1 => n339, IN2 => n338, IN3 => n1131, QN => n341
                           );
   U1062 : OA22X1 port map( IN1 => n1252, IN2 => n1119, IN3 => n1181, IN4 => 
                           n1108, Q => n340);
   U1063 : NAND3X0 port map( IN1 => n341, IN2 => n1128, IN3 => n340, QN => 
                           perm_output(109));
   U1064 : AO22X1 port map( IN1 => eshift_108_port, IN2 => n1031, IN3 => n1020,
                           IN4 => RAMB(97), Q => n342);
   U1065 : AO221X1 port map( IN1 => n1252, IN2 => n1053, IN3 => n1042, IN4 => 
                           RAMB(108), IN5 => n342, Q => n345);
   U1066 : AO22X1 port map( IN1 => addout_108_port, IN2 => n1075, IN3 => 
                           andout_108_port, IN4 => n1064, Q => n343);
   U1067 : AO221X1 port map( IN1 => n213, IN2 => n1097, IN3 => n1086, IN4 => 
                           RAMB(12), IN5 => n343, Q => n344);
   U1068 : OAI21X1 port map( IN1 => n345, IN2 => n344, IN3 => n1131, QN => n347
                           );
   U1069 : OA22X1 port map( IN1 => n1251, IN2 => n1119, IN3 => n1180, IN4 => 
                           n1108, Q => n346);
   U1070 : NAND3X0 port map( IN1 => n347, IN2 => n1128, IN3 => n346, QN => 
                           perm_output(108));
   U1071 : AO22X1 port map( IN1 => eshift_107_port, IN2 => n1031, IN3 => n1020,
                           IN4 => RAMB(96), Q => n348);
   U1072 : AO221X1 port map( IN1 => n1251, IN2 => n1053, IN3 => n1042, IN4 => 
                           RAMB(107), IN5 => n348, Q => n351);
   U1073 : AO22X1 port map( IN1 => addout_107_port, IN2 => n1075, IN3 => 
                           andout_107_port, IN4 => n1064, Q => n349);
   U1074 : AO221X1 port map( IN1 => n87, IN2 => n1097, IN3 => n1086, IN4 => 
                           RAMB(11), IN5 => n349, Q => n350);
   U1075 : OAI21X1 port map( IN1 => n351, IN2 => n350, IN3 => n1132, QN => n353
                           );
   U1076 : OA22X1 port map( IN1 => n1250, IN2 => n1119, IN3 => n1179, IN4 => 
                           n1108, Q => n352);
   U1077 : NAND3X0 port map( IN1 => n353, IN2 => n1128, IN3 => n352, QN => 
                           perm_output(107));
   U1078 : AO22X1 port map( IN1 => eshift_106_port, IN2 => n1031, IN3 => n1020,
                           IN4 => RAMB(127), Q => n354);
   U1079 : AO221X1 port map( IN1 => n1250, IN2 => n1053, IN3 => n1042, IN4 => 
                           RAMB(106), IN5 => n354, Q => n357);
   U1080 : AO22X1 port map( IN1 => addout_106_port, IN2 => n1075, IN3 => 
                           andout_106_port, IN4 => n1064, Q => n355);
   U1081 : AO221X1 port map( IN1 => n106, IN2 => n1097, IN3 => n1086, IN4 => 
                           RAMB(10), IN5 => n355, Q => n356);
   U1082 : OAI21X1 port map( IN1 => n357, IN2 => n356, IN3 => n1132, QN => n359
                           );
   U1083 : OA22X1 port map( IN1 => n1249, IN2 => n1119, IN3 => n1178, IN4 => 
                           n1108, Q => n358);
   U1084 : NAND3X0 port map( IN1 => n359, IN2 => n1128, IN3 => n358, QN => 
                           perm_output(106));
   U1085 : AO22X1 port map( IN1 => eshift_105_port, IN2 => n1031, IN3 => n1020,
                           IN4 => RAMB(126), Q => n360);
   U1086 : AO221X1 port map( IN1 => n1249, IN2 => n1053, IN3 => n1042, IN4 => 
                           RAMB(105), IN5 => n360, Q => n363);
   U1087 : AO22X1 port map( IN1 => n1075, IN2 => addout_105_port, IN3 => 
                           andout_105_port, IN4 => n1064, Q => n361);
   U1088 : AO221X1 port map( IN1 => add_rnd_const_105_port, IN2 => n1097, IN3 
                           => n1086, IN4 => RAMB(9), IN5 => n361, Q => n362);
   U1089 : OAI21X1 port map( IN1 => n363, IN2 => n362, IN3 => n1132, QN => n365
                           );
   U1090 : OA22X1 port map( IN1 => n1248, IN2 => n1119, IN3 => n1177, IN4 => 
                           n1108, Q => n364);
   U1091 : AO22X1 port map( IN1 => eshift_104_port, IN2 => n1031, IN3 => n1020,
                           IN4 => RAMB(125), Q => n366);
   U1092 : AO221X1 port map( IN1 => n1248, IN2 => n1053, IN3 => n1042, IN4 => 
                           RAMB(104), IN5 => n366, Q => n369);
   U1093 : AO22X1 port map( IN1 => addout_104_port, IN2 => n1075, IN3 => 
                           andout_104_port, IN4 => n1064, Q => n367);
   U1094 : AO221X1 port map( IN1 => add_rnd_const_104_port, IN2 => n1097, IN3 
                           => n1086, IN4 => RAMB(8), IN5 => n367, Q => n368);
   U1095 : OAI21X1 port map( IN1 => n369, IN2 => n368, IN3 => n1132, QN => n371
                           );
   U1096 : OA22X1 port map( IN1 => n1247, IN2 => n1119, IN3 => n1176, IN4 => 
                           n1108, Q => n370);
   U1097 : NAND3X0 port map( IN1 => n371, IN2 => n1128, IN3 => n370, QN => 
                           perm_output(104));
   U1098 : AO22X1 port map( IN1 => eshift_103_port, IN2 => n1030, IN3 => n1019,
                           IN4 => RAMB(124), Q => n372);
   U1099 : AO221X1 port map( IN1 => n1247, IN2 => n1052, IN3 => n1041, IN4 => 
                           RAMB(103), IN5 => n372, Q => n375);
   U1100 : AO22X1 port map( IN1 => n1074, IN2 => addout_103_port, IN3 => 
                           andout_103_port, IN4 => n1063, Q => n373);
   U1101 : AO221X1 port map( IN1 => add_rnd_const_103_port, IN2 => n1096, IN3 
                           => n1085, IN4 => RAMB(7), IN5 => n373, Q => n374);
   U1102 : OAI21X1 port map( IN1 => n375, IN2 => n374, IN3 => n1132, QN => n377
                           );
   U1103 : OA22X1 port map( IN1 => n1246, IN2 => n1118, IN3 => n1207, IN4 => 
                           n1107, Q => n376);
   U1104 : NAND3X0 port map( IN1 => n377, IN2 => n1127, IN3 => n376, QN => 
                           perm_output(103));
   U1105 : AO22X1 port map( IN1 => eshift_102_port, IN2 => n1030, IN3 => n1019,
                           IN4 => RAMB(123), Q => n378);
   U1106 : AO221X1 port map( IN1 => n1246, IN2 => n1052, IN3 => n1041, IN4 => 
                           RAMB(102), IN5 => n378, Q => n381);
   U1107 : AO22X1 port map( IN1 => n1074, IN2 => addout_102_port, IN3 => 
                           andout_102_port, IN4 => n1063, Q => n379);
   U1108 : AO221X1 port map( IN1 => add_rnd_const_102_port, IN2 => n1096, IN3 
                           => n1085, IN4 => RAMB(6), IN5 => n379, Q => n380);
   U1109 : OAI21X1 port map( IN1 => n381, IN2 => n380, IN3 => n1132, QN => n383
                           );
   U1110 : OA22X1 port map( IN1 => n1245, IN2 => n1118, IN3 => n1206, IN4 => 
                           n1107, Q => n382);
   U1111 : NAND3X0 port map( IN1 => n383, IN2 => n1127, IN3 => n382, QN => 
                           perm_output(102));
   U1112 : AO22X1 port map( IN1 => eshift_101_port, IN2 => n1030, IN3 => n1019,
                           IN4 => RAMB(122), Q => n384);
   U1113 : AO221X1 port map( IN1 => n1245, IN2 => n1052, IN3 => n1041, IN4 => 
                           RAMB(101), IN5 => n384, Q => n387);
   U1114 : AO22X1 port map( IN1 => addout_101_port, IN2 => n1074, IN3 => 
                           andout_101_port, IN4 => n1063, Q => n385);
   U1115 : AO221X1 port map( IN1 => add_rnd_const_101_port, IN2 => n1096, IN3 
                           => n1085, IN4 => RAMB(5), IN5 => n385, Q => n386);
   U1116 : OAI21X1 port map( IN1 => n387, IN2 => n386, IN3 => n1132, QN => n389
                           );
   U1117 : OA22X1 port map( IN1 => n1244, IN2 => n1118, IN3 => n1205, IN4 => 
                           n1107, Q => n388);
   U1118 : NAND3X0 port map( IN1 => n389, IN2 => n1127, IN3 => n388, QN => 
                           perm_output(101));
   U1119 : AO22X1 port map( IN1 => eshift_100_port, IN2 => n1030, IN3 => n1019,
                           IN4 => RAMB(121), Q => n390);
   U1120 : AO221X1 port map( IN1 => n1244, IN2 => n1052, IN3 => n1041, IN4 => 
                           RAMB(100), IN5 => n390, Q => n393);
   U1121 : AO22X1 port map( IN1 => addout_100_port, IN2 => n1074, IN3 => 
                           andout_100_port, IN4 => n1063, Q => n391);
   U1122 : AO221X1 port map( IN1 => add_rnd_const_100_port, IN2 => n1096, IN3 
                           => n1085, IN4 => RAMB(4), IN5 => n391, Q => n392);
   U1123 : OAI21X1 port map( IN1 => n393, IN2 => n392, IN3 => n1132, QN => n395
                           );
   U1124 : OA22X1 port map( IN1 => n1243, IN2 => n1118, IN3 => n1204, IN4 => 
                           n1107, Q => n394);
   U1125 : NAND3X0 port map( IN1 => n395, IN2 => n1127, IN3 => n394, QN => 
                           perm_output(100));
   U1126 : AO22X1 port map( IN1 => eshift_99_port, IN2 => n1030, IN3 => n1019, 
                           IN4 => RAMB(120), Q => n396);
   U1127 : AO221X1 port map( IN1 => n1243, IN2 => n1052, IN3 => n1041, IN4 => 
                           RAMB(99), IN5 => n396, Q => n399);
   U1128 : AO22X1 port map( IN1 => addout_99_port, IN2 => n1074, IN3 => 
                           andout_99_port, IN4 => n1063, Q => n397);
   U1129 : AO221X1 port map( IN1 => add_rnd_const_99_port, IN2 => n1096, IN3 =>
                           n1085, IN4 => RAMB(3), IN5 => n397, Q => n398);
   U1130 : OAI21X1 port map( IN1 => n399, IN2 => n398, IN3 => n1132, QN => n401
                           );
   U1131 : OA22X1 port map( IN1 => n1242, IN2 => n1118, IN3 => n1203, IN4 => 
                           n1107, Q => n400);
   U1132 : NAND3X0 port map( IN1 => n401, IN2 => n1127, IN3 => n400, QN => 
                           perm_output(99));
   U1133 : AO22X1 port map( IN1 => eshift_98_port, IN2 => n1030, IN3 => n1019, 
                           IN4 => RAMB(119), Q => n402);
   U1134 : AO221X1 port map( IN1 => n1242, IN2 => n1052, IN3 => n1041, IN4 => 
                           RAMB(98), IN5 => n402, Q => n405);
   U1135 : AO22X1 port map( IN1 => addout_98_port, IN2 => n1074, IN3 => 
                           andout_98_port, IN4 => n1063, Q => n403);
   U1136 : AO221X1 port map( IN1 => add_rnd_const_98_port, IN2 => n1096, IN3 =>
                           n1085, IN4 => RAMB(2), IN5 => n403, Q => n404);
   U1137 : OAI21X1 port map( IN1 => n405, IN2 => n404, IN3 => n1132, QN => n407
                           );
   U1138 : OA22X1 port map( IN1 => n1241, IN2 => n1118, IN3 => n1202, IN4 => 
                           n1107, Q => n406);
   U1139 : NAND3X0 port map( IN1 => n407, IN2 => n1127, IN3 => n406, QN => 
                           perm_output(98));
   U1140 : AO22X1 port map( IN1 => eshift_97_port, IN2 => n1030, IN3 => n1019, 
                           IN4 => RAMB(118), Q => n408);
   U1141 : AO221X1 port map( IN1 => n1241, IN2 => n1052, IN3 => n1041, IN4 => 
                           RAMB(97), IN5 => n408, Q => n411);
   U1142 : AO22X1 port map( IN1 => addout_97_port, IN2 => n1074, IN3 => 
                           andout_97_port, IN4 => n1063, Q => n409);
   U1143 : AO221X1 port map( IN1 => add_rnd_const_97_port, IN2 => n1096, IN3 =>
                           n1085, IN4 => RAMB(1), IN5 => n409, Q => n410);
   U1144 : OAI21X1 port map( IN1 => n411, IN2 => n410, IN3 => n1132, QN => n413
                           );
   U1145 : OA22X1 port map( IN1 => n1240, IN2 => n1118, IN3 => n1201, IN4 => 
                           n1107, Q => n412);
   U1146 : NAND3X0 port map( IN1 => n413, IN2 => n1127, IN3 => n412, QN => 
                           perm_output(97));
   U1147 : AO22X1 port map( IN1 => eshift_96_port, IN2 => n1030, IN3 => n1019, 
                           IN4 => RAMB(117), Q => n414);
   U1148 : AO221X1 port map( IN1 => n1240, IN2 => n1052, IN3 => n1041, IN4 => 
                           RAMB(96), IN5 => n414, Q => n417);
   U1149 : AO22X1 port map( IN1 => addout_96_port, IN2 => n1074, IN3 => 
                           andout_96_port, IN4 => n1063, Q => n415);
   U1150 : AO221X1 port map( IN1 => n114, IN2 => n1096, IN3 => n1085, IN4 => 
                           RAMB(0), IN5 => n415, Q => n416);
   U1151 : OAI21X1 port map( IN1 => n417, IN2 => n416, IN3 => n1132, QN => n419
                           );
   U1152 : OA22X1 port map( IN1 => n1271, IN2 => n1118, IN3 => n1200, IN4 => 
                           n1107, Q => n418);
   U1153 : NAND3X0 port map( IN1 => n419, IN2 => n1127, IN3 => n418, QN => 
                           perm_output(96));
   U1154 : AO22X1 port map( IN1 => eshift_95_port, IN2 => n1030, IN3 => n1019, 
                           IN4 => RAMB(84), Q => n420);
   U1155 : AO221X1 port map( IN1 => n1239, IN2 => n1052, IN3 => n1041, IN4 => 
                           RAMB(95), IN5 => n420, Q => n423);
   U1156 : AO22X1 port map( IN1 => addout_95_port, IN2 => n1074, IN3 => 
                           andout_95_port, IN4 => n1063, Q => n421);
   U1157 : AO221X1 port map( IN1 => n212, IN2 => n1096, IN3 => n1085, IN4 => 
                           RAMB(127), IN5 => n421, Q => n422);
   U1158 : OAI21X1 port map( IN1 => n423, IN2 => n422, IN3 => n1133, QN => n425
                           );
   U1159 : OA22X1 port map( IN1 => n1238, IN2 => n1118, IN3 => n1167, IN4 => 
                           n1107, Q => n424);
   U1160 : NAND3X0 port map( IN1 => n425, IN2 => n1127, IN3 => n424, QN => 
                           perm_output(95));
   U1161 : AO22X1 port map( IN1 => eshift_94_port, IN2 => n1030, IN3 => n1019, 
                           IN4 => RAMB(83), Q => n426);
   U1162 : AO221X1 port map( IN1 => n1238, IN2 => n1052, IN3 => n1041, IN4 => 
                           RAMB(94), IN5 => n426, Q => n429);
   U1163 : AO22X1 port map( IN1 => addout_94_port, IN2 => n1074, IN3 => 
                           andout_94_port, IN4 => n1063, Q => n427);
   U1164 : AO221X1 port map( IN1 => n113, IN2 => n1096, IN3 => n1085, IN4 => 
                           RAMB(126), IN5 => n427, Q => n428);
   U1165 : OAI21X1 port map( IN1 => n429, IN2 => n428, IN3 => n1133, QN => n431
                           );
   U1166 : OA22X1 port map( IN1 => n1237, IN2 => n1118, IN3 => n1166, IN4 => 
                           n1107, Q => n430);
   U1167 : NAND3X0 port map( IN1 => n431, IN2 => n1127, IN3 => n430, QN => 
                           perm_output(94));
   U1168 : AO22X1 port map( IN1 => eshift_93_port, IN2 => n1030, IN3 => n1019, 
                           IN4 => RAMB(82), Q => n432);
   U1169 : AO221X1 port map( IN1 => n1237, IN2 => n1052, IN3 => n1041, IN4 => 
                           RAMB(93), IN5 => n432, Q => n435);
   U1170 : AO22X1 port map( IN1 => addout_93_port, IN2 => n1074, IN3 => 
                           andout_93_port, IN4 => n1063, Q => n433);
   U1171 : AO221X1 port map( IN1 => n39, IN2 => n1096, IN3 => n1085, IN4 => 
                           RAMB(125), IN5 => n433, Q => n434);
   U1172 : OAI21X1 port map( IN1 => n435, IN2 => n434, IN3 => n1133, QN => n437
                           );
   U1173 : OA22X1 port map( IN1 => n1236, IN2 => n1118, IN3 => n1165, IN4 => 
                           n1107, Q => n436);
   U1174 : NAND3X0 port map( IN1 => n437, IN2 => n1127, IN3 => n436, QN => 
                           perm_output(93));
   U1175 : AO22X1 port map( IN1 => eshift_92_port, IN2 => n1030, IN3 => n1019, 
                           IN4 => RAMB(81), Q => n438);
   U1176 : AO221X1 port map( IN1 => n1236, IN2 => n1052, IN3 => n1041, IN4 => 
                           RAMB(92), IN5 => n438, Q => n441);
   U1177 : AO22X1 port map( IN1 => addout_92_port, IN2 => n1074, IN3 => 
                           andout_92_port, IN4 => n1063, Q => n439);
   U1178 : AO221X1 port map( IN1 => n218, IN2 => n1096, IN3 => n1085, IN4 => 
                           RAMB(124), IN5 => n439, Q => n440);
   U1179 : OAI21X1 port map( IN1 => n441, IN2 => n440, IN3 => n1133, QN => n443
                           );
   U1180 : OA22X1 port map( IN1 => n1235, IN2 => n1118, IN3 => n1164, IN4 => 
                           n1107, Q => n442);
   U1181 : NAND3X0 port map( IN1 => n443, IN2 => n1127, IN3 => n442, QN => 
                           perm_output(92));
   U1182 : AO22X1 port map( IN1 => eshift_91_port, IN2 => n1029, IN3 => n1018, 
                           IN4 => RAMB(80), Q => n444);
   U1183 : AO221X1 port map( IN1 => n1235, IN2 => n1051, IN3 => n1040, IN4 => 
                           RAMB(91), IN5 => n444, Q => n447);
   U1184 : AO22X1 port map( IN1 => addout_91_port, IN2 => n1073, IN3 => 
                           andout_91_port, IN4 => n1062, Q => n445);
   U1185 : AO221X1 port map( IN1 => n71, IN2 => n1095, IN3 => n1084, IN4 => 
                           RAMB(123), IN5 => n445, Q => n446);
   U1186 : OAI21X1 port map( IN1 => n447, IN2 => n446, IN3 => n1133, QN => n449
                           );
   U1187 : OA22X1 port map( IN1 => n1234, IN2 => n1117, IN3 => n1163, IN4 => 
                           n1106, Q => n448);
   U1188 : NAND3X0 port map( IN1 => n449, IN2 => n1126, IN3 => n448, QN => 
                           perm_output(91));
   U1189 : AO22X1 port map( IN1 => eshift_90_port, IN2 => n1029, IN3 => n1018, 
                           IN4 => RAMB(79), Q => n450);
   U1190 : AO221X1 port map( IN1 => n1234, IN2 => n1051, IN3 => n1040, IN4 => 
                           RAMB(90), IN5 => n450, Q => n453);
   U1191 : AO22X1 port map( IN1 => addout_90_port, IN2 => n1073, IN3 => 
                           andout_90_port, IN4 => n1062, Q => n451);
   U1192 : AO221X1 port map( IN1 => n123, IN2 => n1095, IN3 => n1084, IN4 => 
                           RAMB(122), IN5 => n451, Q => n452);
   U1193 : OAI21X1 port map( IN1 => n453, IN2 => n452, IN3 => n1133, QN => n455
                           );
   U1194 : OA22X1 port map( IN1 => n1233, IN2 => n1117, IN3 => n1162, IN4 => 
                           n1106, Q => n454);
   U1195 : NAND3X0 port map( IN1 => n455, IN2 => n1126, IN3 => n454, QN => 
                           perm_output(90));
   U1196 : AO22X1 port map( IN1 => eshift_89_port, IN2 => n1029, IN3 => n1018, 
                           IN4 => RAMB(78), Q => n456);
   U1197 : AO221X1 port map( IN1 => n1233, IN2 => n1051, IN3 => n1040, IN4 => 
                           RAMB(89), IN5 => n456, Q => n459);
   U1198 : AO22X1 port map( IN1 => addout_89_port, IN2 => n1073, IN3 => 
                           andout_89_port, IN4 => n1062, Q => n457);
   U1199 : AO221X1 port map( IN1 => n66, IN2 => n1095, IN3 => n1084, IN4 => 
                           RAMB(121), IN5 => n457, Q => n458);
   U1200 : OAI21X1 port map( IN1 => n459, IN2 => n458, IN3 => n1133, QN => n461
                           );
   U1201 : OA22X1 port map( IN1 => n1232, IN2 => n1117, IN3 => n1161, IN4 => 
                           n1106, Q => n460);
   U1202 : NAND3X0 port map( IN1 => n461, IN2 => n1126, IN3 => n460, QN => 
                           perm_output(89));
   U1203 : AO22X1 port map( IN1 => eshift_88_port, IN2 => n1029, IN3 => n1018, 
                           IN4 => RAMB(77), Q => n462);
   U1204 : AO221X1 port map( IN1 => n1232, IN2 => n1051, IN3 => n1040, IN4 => 
                           RAMB(88), IN5 => n462, Q => n465);
   U1205 : AO22X1 port map( IN1 => addout_88_port, IN2 => n1073, IN3 => 
                           andout_88_port, IN4 => n1062, Q => n463);
   U1206 : AO221X1 port map( IN1 => n217, IN2 => n1095, IN3 => n1084, IN4 => 
                           RAMB(120), IN5 => n463, Q => n464);
   U1207 : OAI21X1 port map( IN1 => n465, IN2 => n464, IN3 => n1133, QN => n467
                           );
   U1208 : OA22X1 port map( IN1 => n1231, IN2 => n1117, IN3 => n1160, IN4 => 
                           n1106, Q => n466);
   U1209 : AO22X1 port map( IN1 => eshift_87_port, IN2 => n1029, IN3 => n1018, 
                           IN4 => RAMB(76), Q => n468);
   U1210 : AO221X1 port map( IN1 => n1231, IN2 => n1051, IN3 => n1040, IN4 => 
                           RAMB(87), IN5 => n468, Q => n471);
   U1211 : AO22X1 port map( IN1 => addout_87_port, IN2 => n1073, IN3 => 
                           andout_87_port, IN4 => n1062, Q => n469);
   U1212 : AO221X1 port map( IN1 => n77, IN2 => n1095, IN3 => n1084, IN4 => 
                           RAMB(119), IN5 => n469, Q => n470);
   U1213 : OAI21X1 port map( IN1 => n471, IN2 => n470, IN3 => n1133, QN => n473
                           );
   U1214 : OA22X1 port map( IN1 => n1230, IN2 => n1117, IN3 => n1159, IN4 => 
                           n1106, Q => n472);
   U1215 : NAND3X0 port map( IN1 => n473, IN2 => n1126, IN3 => n472, QN => 
                           perm_output(87));
   U1216 : AO22X1 port map( IN1 => eshift_86_port, IN2 => n1029, IN3 => n1018, 
                           IN4 => RAMB(75), Q => n474);
   U1217 : AO221X1 port map( IN1 => n1230, IN2 => n1051, IN3 => n1040, IN4 => 
                           RAMB(86), IN5 => n474, Q => n477);
   U1218 : AO22X1 port map( IN1 => addout_86_port, IN2 => n1073, IN3 => 
                           andout_86_port, IN4 => n1062, Q => n475);
   U1219 : AO221X1 port map( IN1 => n95, IN2 => n1095, IN3 => n1084, IN4 => 
                           RAMB(118), IN5 => n475, Q => n476);
   U1220 : OAI21X1 port map( IN1 => n477, IN2 => n476, IN3 => n1133, QN => n479
                           );
   U1221 : OA22X1 port map( IN1 => n1229, IN2 => n1117, IN3 => n1158, IN4 => 
                           n1106, Q => n478);
   U1222 : NAND3X0 port map( IN1 => n479, IN2 => n1126, IN3 => n478, QN => 
                           perm_output(86));
   U1223 : AO22X1 port map( IN1 => eshift_85_port, IN2 => n1029, IN3 => n1018, 
                           IN4 => RAMB(74), Q => n480);
   U1224 : AO221X1 port map( IN1 => n1229, IN2 => n1051, IN3 => n1040, IN4 => 
                           RAMB(85), IN5 => n480, Q => n483);
   U1225 : AO22X1 port map( IN1 => addout_85_port, IN2 => n1073, IN3 => 
                           andout_85_port, IN4 => n1062, Q => n481);
   U1226 : AO221X1 port map( IN1 => n91, IN2 => n1095, IN3 => n1084, IN4 => 
                           RAMB(117), IN5 => n481, Q => n482);
   U1227 : OAI21X1 port map( IN1 => n483, IN2 => n482, IN3 => n1133, QN => n485
                           );
   U1228 : OA22X1 port map( IN1 => n1228, IN2 => n1117, IN3 => n1157, IN4 => 
                           n1106, Q => n484);
   U1229 : NAND3X0 port map( IN1 => n485, IN2 => n1126, IN3 => n484, QN => 
                           perm_output(85));
   U1230 : AO22X1 port map( IN1 => eshift_84_port, IN2 => n1029, IN3 => n1018, 
                           IN4 => RAMB(73), Q => n486);
   U1231 : AO221X1 port map( IN1 => n1228, IN2 => n1051, IN3 => n1040, IN4 => 
                           RAMB(84), IN5 => n486, Q => n489);
   U1232 : AO22X1 port map( IN1 => addout_84_port, IN2 => n1073, IN3 => 
                           andout_84_port, IN4 => n1062, Q => n487);
   U1233 : AO221X1 port map( IN1 => n33, IN2 => n1095, IN3 => n1084, IN4 => 
                           RAMB(116), IN5 => n487, Q => n488);
   U1234 : OAI21X1 port map( IN1 => n489, IN2 => n488, IN3 => n1133, QN => n491
                           );
   U1235 : OA22X1 port map( IN1 => n1227, IN2 => n1117, IN3 => n1156, IN4 => 
                           n1106, Q => n490);
   U1236 : NAND3X0 port map( IN1 => n491, IN2 => n1126, IN3 => n490, QN => 
                           perm_output(84));
   U1237 : AO22X1 port map( IN1 => eshift_83_port, IN2 => n1029, IN3 => n1018, 
                           IN4 => RAMB(72), Q => n492);
   U1238 : AO221X1 port map( IN1 => n1227, IN2 => n1051, IN3 => n1040, IN4 => 
                           RAMB(83), IN5 => n492, Q => n495);
   U1239 : AO22X1 port map( IN1 => addout_83_port, IN2 => n1073, IN3 => 
                           andout_83_port, IN4 => n1062, Q => n493);
   U1240 : AO221X1 port map( IN1 => n63, IN2 => n1095, IN3 => n1084, IN4 => 
                           RAMB(115), IN5 => n493, Q => n494);
   U1241 : OAI21X1 port map( IN1 => n495, IN2 => n494, IN3 => n1134, QN => n497
                           );
   U1242 : OA22X1 port map( IN1 => n1226, IN2 => n1117, IN3 => n1155, IN4 => 
                           n1106, Q => n496);
   U1243 : NAND3X0 port map( IN1 => n497, IN2 => n1126, IN3 => n496, QN => 
                           perm_output(83));
   U1244 : AO22X1 port map( IN1 => eshift_82_port, IN2 => n1029, IN3 => n1018, 
                           IN4 => RAMB(71), Q => n498);
   U1245 : AO221X1 port map( IN1 => n1226, IN2 => n1051, IN3 => n1040, IN4 => 
                           RAMB(82), IN5 => n498, Q => n501);
   U1246 : AO22X1 port map( IN1 => n1073, IN2 => addout_82_port, IN3 => 
                           andout_82_port, IN4 => n1062, Q => n499);
   U1247 : AO221X1 port map( IN1 => n105, IN2 => n1095, IN3 => n1084, IN4 => 
                           RAMB(114), IN5 => n499, Q => n500);
   U1248 : OAI21X1 port map( IN1 => n501, IN2 => n500, IN3 => n1134, QN => n503
                           );
   U1249 : OA22X1 port map( IN1 => n1225, IN2 => n1117, IN3 => n1154, IN4 => 
                           n1106, Q => n502);
   U1250 : NAND3X0 port map( IN1 => n503, IN2 => n1126, IN3 => n502, QN => 
                           perm_output(82));
   U1251 : AO22X1 port map( IN1 => eshift_81_port, IN2 => n1029, IN3 => n1018, 
                           IN4 => RAMB(70), Q => n504);
   U1252 : AO221X1 port map( IN1 => n1225, IN2 => n1051, IN3 => n1040, IN4 => 
                           RAMB(81), IN5 => n504, Q => n507);
   U1253 : AO22X1 port map( IN1 => addout_81_port, IN2 => n1073, IN3 => 
                           andout_81_port, IN4 => n1062, Q => n505);
   U1254 : AO221X1 port map( IN1 => n118, IN2 => n1095, IN3 => n1084, IN4 => 
                           RAMB(113), IN5 => n505, Q => n506);
   U1255 : OAI21X1 port map( IN1 => n507, IN2 => n506, IN3 => n1134, QN => n509
                           );
   U1256 : OA22X1 port map( IN1 => n1224, IN2 => n1117, IN3 => n1153, IN4 => 
                           n1106, Q => n508);
   U1257 : NAND3X0 port map( IN1 => n509, IN2 => n1126, IN3 => n508, QN => 
                           perm_output(81));
   U1258 : AO22X1 port map( IN1 => eshift_80_port, IN2 => n1029, IN3 => n1018, 
                           IN4 => RAMB(69), Q => n510);
   U1259 : AO221X1 port map( IN1 => n1224, IN2 => n1051, IN3 => n1040, IN4 => 
                           RAMB(80), IN5 => n510, Q => n513);
   U1260 : AO22X1 port map( IN1 => addout_80_port, IN2 => n1073, IN3 => 
                           andout_80_port, IN4 => n1062, Q => n511);
   U1261 : AO221X1 port map( IN1 => n56, IN2 => n1095, IN3 => n1084, IN4 => 
                           RAMB(112), IN5 => n511, Q => n512);
   U1262 : OAI21X1 port map( IN1 => n513, IN2 => n512, IN3 => n1134, QN => n515
                           );
   U1263 : OA22X1 port map( IN1 => n1223, IN2 => n1117, IN3 => n1152, IN4 => 
                           n1106, Q => n514);
   U1264 : NAND3X0 port map( IN1 => n515, IN2 => n1126, IN3 => n514, QN => 
                           perm_output(80));
   U1265 : AO22X1 port map( IN1 => eshift_79_port, IN2 => n1028, IN3 => n1017, 
                           IN4 => RAMB(68), Q => n516);
   U1266 : AO221X1 port map( IN1 => n1223, IN2 => n1050, IN3 => n1039, IN4 => 
                           RAMB(79), IN5 => n516, Q => n519);
   U1267 : AO22X1 port map( IN1 => addout_79_port, IN2 => n1072, IN3 => 
                           andout_79_port, IN4 => n1061, Q => n517);
   U1268 : AO221X1 port map( IN1 => n115, IN2 => n1094, IN3 => n1083, IN4 => 
                           RAMB(111), IN5 => n517, Q => n518);
   U1269 : OAI21X1 port map( IN1 => n519, IN2 => n518, IN3 => n1134, QN => n521
                           );
   U1270 : OA22X1 port map( IN1 => n1222, IN2 => n1116, IN3 => n1151, IN4 => 
                           n1105, Q => n520);
   U1271 : NAND3X0 port map( IN1 => n521, IN2 => n1125, IN3 => n520, QN => 
                           perm_output(79));
   U1272 : AO22X1 port map( IN1 => eshift_78_port, IN2 => n1028, IN3 => n1017, 
                           IN4 => RAMB(67), Q => n522);
   U1273 : AO221X1 port map( IN1 => n1222, IN2 => n1050, IN3 => n1039, IN4 => 
                           RAMB(78), IN5 => n522, Q => n525);
   U1274 : AO22X1 port map( IN1 => addout_78_port, IN2 => n1072, IN3 => 
                           andout_78_port, IN4 => n1061, Q => n523);
   U1275 : AO221X1 port map( IN1 => n107, IN2 => n1094, IN3 => n1083, IN4 => 
                           RAMB(110), IN5 => n523, Q => n524);
   U1276 : OAI21X1 port map( IN1 => n525, IN2 => n524, IN3 => n1134, QN => n527
                           );
   U1277 : OA22X1 port map( IN1 => n1221, IN2 => n1116, IN3 => n1150, IN4 => 
                           n1105, Q => n526);
   U1278 : NAND3X0 port map( IN1 => n527, IN2 => n1125, IN3 => n526, QN => 
                           perm_output(78));
   U1279 : AO22X1 port map( IN1 => eshift_77_port, IN2 => n1028, IN3 => n1017, 
                           IN4 => RAMB(66), Q => n528);
   U1280 : AO221X1 port map( IN1 => n1221, IN2 => n1050, IN3 => n1039, IN4 => 
                           RAMB(77), IN5 => n528, Q => n531);
   U1281 : AO22X1 port map( IN1 => addout_77_port, IN2 => n1072, IN3 => 
                           andout_77_port, IN4 => n1061, Q => n529);
   U1282 : AO221X1 port map( IN1 => n62, IN2 => n1094, IN3 => n1083, IN4 => 
                           RAMB(109), IN5 => n529, Q => n530);
   U1283 : OAI21X1 port map( IN1 => n531, IN2 => n530, IN3 => n1134, QN => n533
                           );
   U1284 : OA22X1 port map( IN1 => n1220, IN2 => n1116, IN3 => n1149, IN4 => 
                           n1105, Q => n532);
   U1285 : NAND3X0 port map( IN1 => n533, IN2 => n1125, IN3 => n532, QN => 
                           perm_output(77));
   U1286 : AO22X1 port map( IN1 => eshift_76_port, IN2 => n1028, IN3 => n1017, 
                           IN4 => RAMB(65), Q => n534);
   U1287 : AO221X1 port map( IN1 => n1220, IN2 => n1050, IN3 => n1039, IN4 => 
                           RAMB(76), IN5 => n534, Q => n537);
   U1288 : AO22X1 port map( IN1 => addout_76_port, IN2 => n1072, IN3 => 
                           andout_76_port, IN4 => n1061, Q => n535);
   U1289 : AO221X1 port map( IN1 => n137, IN2 => n1094, IN3 => n1083, IN4 => 
                           RAMB(108), IN5 => n535, Q => n536);
   U1290 : OAI21X1 port map( IN1 => n537, IN2 => n536, IN3 => n1134, QN => n539
                           );
   U1291 : OA22X1 port map( IN1 => n1219, IN2 => n1116, IN3 => n1148, IN4 => 
                           n1105, Q => n538);
   U1292 : NAND3X0 port map( IN1 => n539, IN2 => n1125, IN3 => n538, QN => 
                           perm_output(76));
   U1293 : AO22X1 port map( IN1 => eshift_75_port, IN2 => n1028, IN3 => n1017, 
                           IN4 => RAMB(64), Q => n540);
   U1294 : AO221X1 port map( IN1 => n1219, IN2 => n1050, IN3 => n1039, IN4 => 
                           RAMB(75), IN5 => n540, Q => n543);
   U1295 : AO22X1 port map( IN1 => addout_75_port, IN2 => n1072, IN3 => 
                           andout_75_port, IN4 => n1061, Q => n541);
   U1296 : AO221X1 port map( IN1 => n42, IN2 => n1094, IN3 => n1083, IN4 => 
                           RAMB(107), IN5 => n541, Q => n542);
   U1297 : OAI21X1 port map( IN1 => n543, IN2 => n542, IN3 => n1134, QN => n545
                           );
   U1298 : OA22X1 port map( IN1 => n1218, IN2 => n1116, IN3 => n1147, IN4 => 
                           n1105, Q => n544);
   U1299 : AO22X1 port map( IN1 => eshift_74_port, IN2 => n1028, IN3 => n1017, 
                           IN4 => RAMB(95), Q => n546);
   U1300 : AO221X1 port map( IN1 => n1218, IN2 => n1050, IN3 => n1039, IN4 => 
                           RAMB(74), IN5 => n546, Q => n549);
   U1301 : AO22X1 port map( IN1 => addout_74_port, IN2 => n1072, IN3 => 
                           andout_74_port, IN4 => n1061, Q => n547);
   U1302 : AO221X1 port map( IN1 => n139, IN2 => n1094, IN3 => n1083, IN4 => 
                           RAMB(106), IN5 => n547, Q => n548);
   U1303 : OAI21X1 port map( IN1 => n549, IN2 => n548, IN3 => n1134, QN => n551
                           );
   U1304 : OA22X1 port map( IN1 => n1217, IN2 => n1116, IN3 => n1146, IN4 => 
                           n1105, Q => n550);
   U1305 : NAND3X0 port map( IN1 => n551, IN2 => n1125, IN3 => n550, QN => 
                           perm_output(74));
   U1306 : AO22X1 port map( IN1 => eshift_73_port, IN2 => n1028, IN3 => n1017, 
                           IN4 => RAMB(94), Q => n552);
   U1307 : AO221X1 port map( IN1 => n1217, IN2 => n1050, IN3 => n1039, IN4 => 
                           RAMB(73), IN5 => n552, Q => n555);
   U1308 : AO22X1 port map( IN1 => addout_73_port, IN2 => n1072, IN3 => 
                           andout_73_port, IN4 => n1061, Q => n553);
   U1309 : AO221X1 port map( IN1 => n110, IN2 => n1094, IN3 => n1083, IN4 => 
                           RAMB(105), IN5 => n553, Q => n554);
   U1310 : OAI21X1 port map( IN1 => n555, IN2 => n554, IN3 => n1134, QN => n557
                           );
   U1311 : OA22X1 port map( IN1 => n1216, IN2 => n1116, IN3 => n1145, IN4 => 
                           n1105, Q => n556);
   U1312 : NAND3X0 port map( IN1 => n557, IN2 => n1125, IN3 => n556, QN => 
                           perm_output(73));
   U1313 : AO22X1 port map( IN1 => eshift_72_port, IN2 => n1028, IN3 => n1017, 
                           IN4 => RAMB(93), Q => n558);
   U1314 : AO221X1 port map( IN1 => n1216, IN2 => n1050, IN3 => n1039, IN4 => 
                           RAMB(72), IN5 => n558, Q => n561);
   U1315 : AO22X1 port map( IN1 => addout_72_port, IN2 => n1072, IN3 => 
                           andout_72_port, IN4 => n1061, Q => n559);
   U1316 : AO221X1 port map( IN1 => n128, IN2 => n1094, IN3 => n1083, IN4 => 
                           RAMB(104), IN5 => n559, Q => n560);
   U1317 : OAI21X1 port map( IN1 => n561, IN2 => n560, IN3 => n1134, QN => n563
                           );
   U1318 : OA22X1 port map( IN1 => n1215, IN2 => n1116, IN3 => n1144, IN4 => 
                           n1105, Q => n562);
   U1319 : NAND3X0 port map( IN1 => n563, IN2 => n1125, IN3 => n562, QN => 
                           perm_output(72));
   U1320 : AO22X1 port map( IN1 => eshift_71_port, IN2 => n1028, IN3 => n1017, 
                           IN4 => RAMB(92), Q => n564);
   U1321 : AO221X1 port map( IN1 => n1215, IN2 => n1050, IN3 => n1039, IN4 => 
                           RAMB(71), IN5 => n564, Q => n567);
   U1322 : AO22X1 port map( IN1 => addout_71_port, IN2 => n1072, IN3 => 
                           andout_71_port, IN4 => n1061, Q => n565);
   U1323 : AO221X1 port map( IN1 => n19, IN2 => n1094, IN3 => n1083, IN4 => 
                           RAMB(103), IN5 => n565, Q => n566);
   U1324 : OAI21X1 port map( IN1 => n567, IN2 => n566, IN3 => n1135, QN => n569
                           );
   U1325 : OA22X1 port map( IN1 => n1214, IN2 => n1116, IN3 => n1175, IN4 => 
                           n1105, Q => n568);
   U1326 : NAND3X0 port map( IN1 => n569, IN2 => n1125, IN3 => n568, QN => 
                           perm_output(71));
   U1327 : AO22X1 port map( IN1 => eshift_70_port, IN2 => n1028, IN3 => n1017, 
                           IN4 => RAMB(91), Q => n570);
   U1328 : AO221X1 port map( IN1 => n1214, IN2 => n1050, IN3 => n1039, IN4 => 
                           RAMB(70), IN5 => n570, Q => n573);
   U1329 : AO22X1 port map( IN1 => addout_70_port, IN2 => n1072, IN3 => 
                           andout_70_port, IN4 => n1061, Q => n571);
   U1330 : AO221X1 port map( IN1 => n58, IN2 => n1094, IN3 => n1083, IN4 => 
                           RAMB(102), IN5 => n571, Q => n572);
   U1331 : OAI21X1 port map( IN1 => n573, IN2 => n572, IN3 => n1135, QN => n575
                           );
   U1332 : OA22X1 port map( IN1 => n1213, IN2 => n1116, IN3 => n1174, IN4 => 
                           n1105, Q => n574);
   U1333 : NAND3X0 port map( IN1 => n575, IN2 => n1125, IN3 => n574, QN => 
                           perm_output(70));
   U1334 : AO22X1 port map( IN1 => eshift_69_port, IN2 => n1028, IN3 => n1017, 
                           IN4 => RAMB(90), Q => n576);
   U1335 : AO221X1 port map( IN1 => n1213, IN2 => n1050, IN3 => n1039, IN4 => 
                           RAMB(69), IN5 => n576, Q => n579);
   U1336 : AO22X1 port map( IN1 => addout_69_port, IN2 => n1072, IN3 => 
                           andout_69_port, IN4 => n1061, Q => n577);
   U1337 : AO221X1 port map( IN1 => n109, IN2 => n1094, IN3 => n1083, IN4 => 
                           RAMB(101), IN5 => n577, Q => n578);
   U1338 : OAI21X1 port map( IN1 => n579, IN2 => n578, IN3 => n1135, QN => n581
                           );
   U1339 : OA22X1 port map( IN1 => n1212, IN2 => n1116, IN3 => n1173, IN4 => 
                           n1105, Q => n580);
   U1340 : NAND3X0 port map( IN1 => n581, IN2 => n1125, IN3 => n580, QN => 
                           perm_output(69));
   U1341 : AO22X1 port map( IN1 => eshift_68_port, IN2 => n1028, IN3 => n1017, 
                           IN4 => RAMB(89), Q => n582);
   U1342 : AO221X1 port map( IN1 => n1212, IN2 => n1050, IN3 => n1039, IN4 => 
                           RAMB(68), IN5 => n582, Q => n585);
   U1343 : AO22X1 port map( IN1 => addout_68_port, IN2 => n1072, IN3 => 
                           andout_68_port, IN4 => n1061, Q => n583);
   U1344 : AO221X1 port map( IN1 => n220, IN2 => n1094, IN3 => n1083, IN4 => 
                           RAMB(100), IN5 => n583, Q => n584);
   U1345 : OAI21X1 port map( IN1 => n585, IN2 => n584, IN3 => n1135, QN => n587
                           );
   U1346 : OA22X1 port map( IN1 => n1211, IN2 => n1116, IN3 => n1172, IN4 => 
                           n1105, Q => n586);
   U1347 : NAND3X0 port map( IN1 => n587, IN2 => n1125, IN3 => n586, QN => 
                           perm_output(68));
   U1348 : AO22X1 port map( IN1 => eshift_67_port, IN2 => n1027, IN3 => n1016, 
                           IN4 => RAMB(88), Q => n588);
   U1349 : AO221X1 port map( IN1 => n1211, IN2 => n1049, IN3 => n1038, IN4 => 
                           RAMB(67), IN5 => n588, Q => n591);
   U1350 : AO22X1 port map( IN1 => addout_67_port, IN2 => n1071, IN3 => 
                           andout_67_port, IN4 => n1060, Q => n589);
   U1351 : AO221X1 port map( IN1 => n79, IN2 => n1093, IN3 => n1082, IN4 => 
                           RAMB(99), IN5 => n589, Q => n590);
   U1352 : OAI21X1 port map( IN1 => n591, IN2 => n590, IN3 => n1135, QN => n593
                           );
   U1353 : OA22X1 port map( IN1 => n1210, IN2 => n1115, IN3 => n1171, IN4 => 
                           n1104, Q => n592);
   U1354 : NAND3X0 port map( IN1 => n593, IN2 => n1124, IN3 => n592, QN => 
                           perm_output(67));
   U1355 : AO22X1 port map( IN1 => eshift_66_port, IN2 => n1027, IN3 => n1016, 
                           IN4 => RAMB(87), Q => n594);
   U1356 : AO221X1 port map( IN1 => n1210, IN2 => n1049, IN3 => n1038, IN4 => 
                           RAMB(66), IN5 => n594, Q => n597);
   U1357 : AO22X1 port map( IN1 => addout_66_port, IN2 => n1071, IN3 => 
                           andout_66_port, IN4 => n1060, Q => n595);
   U1358 : AO221X1 port map( IN1 => n223, IN2 => n1093, IN3 => n1082, IN4 => 
                           RAMB(98), IN5 => n595, Q => n596);
   U1359 : OAI21X1 port map( IN1 => n597, IN2 => n596, IN3 => n1135, QN => n599
                           );
   U1360 : OA22X1 port map( IN1 => n1209, IN2 => n1115, IN3 => n1170, IN4 => 
                           n1104, Q => n598);
   U1361 : NAND3X0 port map( IN1 => n599, IN2 => n1124, IN3 => n598, QN => 
                           perm_output(66));
   U1362 : AO22X1 port map( IN1 => eshift_65_port, IN2 => n1027, IN3 => n1016, 
                           IN4 => RAMB(86), Q => n600);
   U1363 : AO221X1 port map( IN1 => n1209, IN2 => n1049, IN3 => n1038, IN4 => 
                           RAMB(65), IN5 => n600, Q => n603);
   U1364 : AO22X1 port map( IN1 => addout_65_port, IN2 => n1071, IN3 => 
                           andout_65_port, IN4 => n1060, Q => n601);
   U1365 : AO221X1 port map( IN1 => n49, IN2 => n1093, IN3 => n1082, IN4 => 
                           RAMB(97), IN5 => n601, Q => n602);
   U1366 : OAI21X1 port map( IN1 => n603, IN2 => n602, IN3 => n1135, QN => n605
                           );
   U1367 : OA22X1 port map( IN1 => n1208, IN2 => n1115, IN3 => n1169, IN4 => 
                           n1104, Q => n604);
   U1368 : NAND3X0 port map( IN1 => n605, IN2 => n1124, IN3 => n604, QN => 
                           perm_output(65));
   U1369 : AO22X1 port map( IN1 => eshift_64_port, IN2 => n1027, IN3 => n1016, 
                           IN4 => RAMB(85), Q => n606);
   U1370 : AO221X1 port map( IN1 => n1208, IN2 => n1049, IN3 => n1038, IN4 => 
                           RAMB(64), IN5 => n606, Q => n609);
   U1371 : AO22X1 port map( IN1 => addout_64_port, IN2 => n1071, IN3 => 
                           andout_64_port, IN4 => n1060, Q => n607);
   U1372 : AO221X1 port map( IN1 => n121, IN2 => n1093, IN3 => n1082, IN4 => 
                           RAMB(96), IN5 => n607, Q => n608);
   U1373 : OAI21X1 port map( IN1 => n609, IN2 => n608, IN3 => n1135, QN => n611
                           );
   U1374 : OA22X1 port map( IN1 => n1239, IN2 => n1115, IN3 => n1168, IN4 => 
                           n1104, Q => n610);
   U1375 : NAND3X0 port map( IN1 => n611, IN2 => n1124, IN3 => n610, QN => 
                           perm_output(64));
   U1376 : AO22X1 port map( IN1 => eshift_63_port, IN2 => n1027, IN3 => n1016, 
                           IN4 => RAMB(52), Q => n612);
   U1377 : AO221X1 port map( IN1 => n1207, IN2 => n1049, IN3 => n1038, IN4 => 
                           RAMB(63), IN5 => n612, Q => n615);
   U1378 : AO22X1 port map( IN1 => addout_63_port, IN2 => n1071, IN3 => 
                           andout_63_port, IN4 => n1060, Q => n613);
   U1379 : AO221X1 port map( IN1 => n78, IN2 => n1093, IN3 => n1082, IN4 => 
                           RAMB(95), IN5 => n613, Q => n614);
   U1380 : OAI21X1 port map( IN1 => n615, IN2 => n614, IN3 => n1135, QN => n617
                           );
   U1381 : OA22X1 port map( IN1 => n1206, IN2 => n1115, IN3 => n1263, IN4 => 
                           n1104, Q => n616);
   U1382 : NAND3X0 port map( IN1 => n617, IN2 => n1124, IN3 => n616, QN => 
                           perm_output(63));
   U1383 : AO22X1 port map( IN1 => eshift_62_port, IN2 => n1027, IN3 => n1016, 
                           IN4 => RAMB(51), Q => n618);
   U1384 : AO221X1 port map( IN1 => n1206, IN2 => n1049, IN3 => n1038, IN4 => 
                           RAMB(62), IN5 => n618, Q => n621);
   U1385 : AO22X1 port map( IN1 => addout_62_port, IN2 => n1071, IN3 => 
                           andout_62_port, IN4 => n1060, Q => n619);
   U1386 : AO221X1 port map( IN1 => n52, IN2 => n1093, IN3 => n1082, IN4 => 
                           RAMB(94), IN5 => n619, Q => n620);
   U1387 : OAI21X1 port map( IN1 => n621, IN2 => n620, IN3 => n1135, QN => n623
                           );
   U1388 : OA22X1 port map( IN1 => n1205, IN2 => n1115, IN3 => n1262, IN4 => 
                           n1104, Q => n622);
   U1389 : NAND3X0 port map( IN1 => n623, IN2 => n1124, IN3 => n622, QN => 
                           perm_output(62));
   U1390 : AO22X1 port map( IN1 => eshift_61_port, IN2 => n1027, IN3 => n1016, 
                           IN4 => RAMB(50), Q => n624);
   U1391 : AO221X1 port map( IN1 => n1205, IN2 => n1049, IN3 => n1038, IN4 => 
                           RAMB(61), IN5 => n624, Q => n627);
   U1392 : AO22X1 port map( IN1 => addout_61_port, IN2 => n1071, IN3 => 
                           andout_61_port, IN4 => n1060, Q => n625);
   U1393 : AO221X1 port map( IN1 => n100, IN2 => n1093, IN3 => n1082, IN4 => 
                           RAMB(93), IN5 => n625, Q => n626);
   U1394 : OAI21X1 port map( IN1 => n627, IN2 => n626, IN3 => n1135, QN => n629
                           );
   U1395 : OA22X1 port map( IN1 => n1204, IN2 => n1115, IN3 => n1261, IN4 => 
                           n1104, Q => n628);
   U1396 : NAND3X0 port map( IN1 => n629, IN2 => n1124, IN3 => n628, QN => 
                           perm_output(61));
   U1397 : AO22X1 port map( IN1 => eshift_60_port, IN2 => n1027, IN3 => n1016, 
                           IN4 => RAMB(49), Q => n630);
   U1398 : AO221X1 port map( IN1 => n1204, IN2 => n1049, IN3 => n1038, IN4 => 
                           RAMB(60), IN5 => n630, Q => n633);
   U1399 : AO22X1 port map( IN1 => addout_60_port, IN2 => n1071, IN3 => 
                           andout_60_port, IN4 => n1060, Q => n631);
   U1400 : AO221X1 port map( IN1 => n81, IN2 => n1093, IN3 => n1082, IN4 => 
                           RAMB(92), IN5 => n631, Q => n632);
   U1401 : OAI21X1 port map( IN1 => n633, IN2 => n632, IN3 => n1135, QN => n635
                           );
   U1402 : OA22X1 port map( IN1 => n1203, IN2 => n1115, IN3 => n1260, IN4 => 
                           n1104, Q => n634);
   U1403 : NAND3X0 port map( IN1 => n635, IN2 => n1124, IN3 => n634, QN => 
                           perm_output(60));
   U1404 : AO22X1 port map( IN1 => eshift_59_port, IN2 => n1027, IN3 => n1016, 
                           IN4 => RAMB(48), Q => n636);
   U1405 : AO221X1 port map( IN1 => n1203, IN2 => n1049, IN3 => n1038, IN4 => 
                           RAMB(59), IN5 => n636, Q => n639);
   U1406 : AO22X1 port map( IN1 => addout_59_port, IN2 => n1071, IN3 => 
                           andout_59_port, IN4 => n1060, Q => n637);
   U1407 : AO221X1 port map( IN1 => n53, IN2 => n1093, IN3 => n1082, IN4 => 
                           RAMB(91), IN5 => n637, Q => n638);
   U1408 : OAI21X1 port map( IN1 => n639, IN2 => n638, IN3 => n1136, QN => n641
                           );
   U1409 : OA22X1 port map( IN1 => n1202, IN2 => n1115, IN3 => n1259, IN4 => 
                           n1104, Q => n640);
   U1410 : NAND3X0 port map( IN1 => n641, IN2 => n1124, IN3 => n640, QN => 
                           perm_output(59));
   U1411 : AO22X1 port map( IN1 => eshift_58_port, IN2 => n1027, IN3 => n1016, 
                           IN4 => RAMB(47), Q => n642);
   U1412 : AO221X1 port map( IN1 => n1202, IN2 => n1049, IN3 => n1038, IN4 => 
                           RAMB(58), IN5 => n642, Q => n645);
   U1413 : AO22X1 port map( IN1 => addout_58_port, IN2 => n1071, IN3 => 
                           andout_58_port, IN4 => n1060, Q => n643);
   U1414 : AO221X1 port map( IN1 => n124, IN2 => n1093, IN3 => n1082, IN4 => 
                           RAMB(90), IN5 => n643, Q => n644);
   U1415 : OAI21X1 port map( IN1 => n645, IN2 => n644, IN3 => n1136, QN => n647
                           );
   U1416 : OA22X1 port map( IN1 => n1201, IN2 => n1115, IN3 => n1258, IN4 => 
                           n1104, Q => n646);
   U1417 : NAND3X0 port map( IN1 => n647, IN2 => n1124, IN3 => n646, QN => 
                           perm_output(58));
   U1418 : AO22X1 port map( IN1 => eshift_57_port, IN2 => n1027, IN3 => n1016, 
                           IN4 => RAMB(46), Q => n648);
   U1419 : AO221X1 port map( IN1 => n1201, IN2 => n1049, IN3 => n1038, IN4 => 
                           RAMB(57), IN5 => n648, Q => n651);
   U1420 : AO22X1 port map( IN1 => n1071, IN2 => addout_57_port, IN3 => 
                           andout_57_port, IN4 => n1060, Q => n649);
   U1421 : AO221X1 port map( IN1 => n207, IN2 => n1093, IN3 => n1082, IN4 => 
                           RAMB(89), IN5 => n649, Q => n650);
   U1422 : OAI21X1 port map( IN1 => n651, IN2 => n650, IN3 => n1136, QN => n653
                           );
   U1423 : OA22X1 port map( IN1 => n1200, IN2 => n1115, IN3 => n1257, IN4 => 
                           n1104, Q => n652);
   U1424 : AO22X1 port map( IN1 => eshift_56_port, IN2 => n1027, IN3 => n1016, 
                           IN4 => RAMB(45), Q => n654);
   U1425 : AO221X1 port map( IN1 => n1200, IN2 => n1049, IN3 => n1038, IN4 => 
                           RAMB(56), IN5 => n654, Q => n657);
   U1426 : AO22X1 port map( IN1 => addout_56_port, IN2 => n1071, IN3 => 
                           andout_56_port, IN4 => n1060, Q => n655);
   U1427 : AO221X1 port map( IN1 => n136, IN2 => n1093, IN3 => n1082, IN4 => 
                           RAMB(88), IN5 => n655, Q => n656);
   U1428 : OAI21X1 port map( IN1 => n657, IN2 => n656, IN3 => n1136, QN => n659
                           );
   U1429 : OA22X1 port map( IN1 => n1199, IN2 => n1115, IN3 => n1256, IN4 => 
                           n1104, Q => n658);
   U1430 : NAND3X0 port map( IN1 => n659, IN2 => n1124, IN3 => n658, QN => 
                           perm_output(56));
   U1431 : AO22X1 port map( IN1 => eshift_55_port, IN2 => n1026, IN3 => n1015, 
                           IN4 => RAMB(44), Q => n660);
   U1432 : AO221X1 port map( IN1 => n1199, IN2 => n1048, IN3 => n1037, IN4 => 
                           RAMB(55), IN5 => n660, Q => n663);
   U1433 : AO22X1 port map( IN1 => addout_55_port, IN2 => n1070, IN3 => 
                           andout_55_port, IN4 => n1059, Q => n661);
   U1434 : AO221X1 port map( IN1 => n69, IN2 => n1092, IN3 => n1081, IN4 => 
                           RAMB(87), IN5 => n661, Q => n662);
   U1435 : OAI21X1 port map( IN1 => n663, IN2 => n662, IN3 => n1136, QN => n665
                           );
   U1436 : OA22X1 port map( IN1 => n1198, IN2 => n1114, IN3 => n1255, IN4 => 
                           n1103, Q => n664);
   U1437 : NAND3X0 port map( IN1 => n665, IN2 => n1123, IN3 => n664, QN => 
                           perm_output(55));
   U1438 : AO22X1 port map( IN1 => eshift_54_port, IN2 => n1026, IN3 => n1015, 
                           IN4 => RAMB(43), Q => n666);
   U1439 : AO221X1 port map( IN1 => n1198, IN2 => n1048, IN3 => n1037, IN4 => 
                           RAMB(54), IN5 => n666, Q => n669);
   U1440 : AO22X1 port map( IN1 => addout_54_port, IN2 => n1070, IN3 => 
                           andout_54_port, IN4 => n1059, Q => n667);
   U1441 : AO221X1 port map( IN1 => n54, IN2 => n1092, IN3 => n1081, IN4 => 
                           RAMB(86), IN5 => n667, Q => n668);
   U1442 : OAI21X1 port map( IN1 => n669, IN2 => n668, IN3 => n1136, QN => n671
                           );
   U1443 : OA22X1 port map( IN1 => n1197, IN2 => n1114, IN3 => n1254, IN4 => 
                           n1103, Q => n670);
   U1444 : NAND3X0 port map( IN1 => n671, IN2 => n1123, IN3 => n670, QN => 
                           perm_output(54));
   U1445 : AO22X1 port map( IN1 => eshift_53_port, IN2 => n1026, IN3 => n1015, 
                           IN4 => RAMB(42), Q => n672);
   U1446 : AO221X1 port map( IN1 => n1197, IN2 => n1048, IN3 => n1037, IN4 => 
                           RAMB(53), IN5 => n672, Q => n675);
   U1447 : AO22X1 port map( IN1 => addout_53_port, IN2 => n1070, IN3 => 
                           andout_53_port, IN4 => n1059, Q => n673);
   U1448 : AO221X1 port map( IN1 => n131, IN2 => n1092, IN3 => n1081, IN4 => 
                           RAMB(85), IN5 => n673, Q => n674);
   U1449 : OAI21X1 port map( IN1 => n675, IN2 => n674, IN3 => n1136, QN => n677
                           );
   U1450 : OA22X1 port map( IN1 => n1196, IN2 => n1114, IN3 => n1253, IN4 => 
                           n1103, Q => n676);
   U1451 : NAND3X0 port map( IN1 => n677, IN2 => n1123, IN3 => n676, QN => 
                           perm_output(53));
   U1452 : AO22X1 port map( IN1 => eshift_52_port, IN2 => n1026, IN3 => n1015, 
                           IN4 => RAMB(41), Q => n678);
   U1453 : AO221X1 port map( IN1 => n1196, IN2 => n1048, IN3 => n1037, IN4 => 
                           RAMB(52), IN5 => n678, Q => n681);
   U1454 : AO22X1 port map( IN1 => addout_52_port, IN2 => n1070, IN3 => 
                           andout_52_port, IN4 => n1059, Q => n679);
   U1455 : AO221X1 port map( IN1 => n31, IN2 => n1092, IN3 => n1081, IN4 => 
                           RAMB(84), IN5 => n679, Q => n680);
   U1456 : OAI21X1 port map( IN1 => n681, IN2 => n680, IN3 => n1136, QN => n683
                           );
   U1457 : OA22X1 port map( IN1 => n1195, IN2 => n1114, IN3 => n1252, IN4 => 
                           n1103, Q => n682);
   U1458 : NAND3X0 port map( IN1 => n683, IN2 => n1123, IN3 => n682, QN => 
                           perm_output(52));
   U1459 : AO22X1 port map( IN1 => eshift_51_port, IN2 => n1026, IN3 => n1015, 
                           IN4 => RAMB(40), Q => n684);
   U1460 : AO221X1 port map( IN1 => n1195, IN2 => n1048, IN3 => n1037, IN4 => 
                           RAMB(51), IN5 => n684, Q => n687);
   U1461 : AO22X1 port map( IN1 => addout_51_port, IN2 => n1070, IN3 => 
                           andout_51_port, IN4 => n1059, Q => n685);
   U1462 : AO221X1 port map( IN1 => n133, IN2 => n1092, IN3 => n1081, IN4 => 
                           RAMB(83), IN5 => n685, Q => n686);
   U1463 : OAI21X1 port map( IN1 => n687, IN2 => n686, IN3 => n1136, QN => n689
                           );
   U1464 : OA22X1 port map( IN1 => n1194, IN2 => n1114, IN3 => n1251, IN4 => 
                           n1103, Q => n688);
   U1465 : NAND3X0 port map( IN1 => n689, IN2 => n1123, IN3 => n688, QN => 
                           perm_output(51));
   U1466 : AO22X1 port map( IN1 => eshift_50_port, IN2 => n1026, IN3 => n1015, 
                           IN4 => n16, Q => n690);
   U1467 : AO221X1 port map( IN1 => n1194, IN2 => n1048, IN3 => n1037, IN4 => 
                           RAMB(50), IN5 => n690, Q => n693);
   U1468 : AO22X1 port map( IN1 => addout_50_port, IN2 => n1070, IN3 => 
                           andout_50_port, IN4 => n1059, Q => n691);
   U1469 : AO221X1 port map( IN1 => n116, IN2 => n1092, IN3 => n1081, IN4 => 
                           RAMB(82), IN5 => n691, Q => n692);
   U1470 : OAI21X1 port map( IN1 => n693, IN2 => n692, IN3 => n1136, QN => n695
                           );
   U1471 : OA22X1 port map( IN1 => n1193, IN2 => n1114, IN3 => n1250, IN4 => 
                           n1103, Q => n694);
   U1472 : NAND3X0 port map( IN1 => n695, IN2 => n1123, IN3 => n694, QN => 
                           perm_output(50));
   U1473 : AO22X1 port map( IN1 => eshift_49_port, IN2 => n1026, IN3 => n1015, 
                           IN4 => RAMB(38), Q => n696);
   U1474 : AO221X1 port map( IN1 => n1193, IN2 => n1048, IN3 => n1037, IN4 => 
                           RAMB(49), IN5 => n696, Q => n699);
   U1475 : AO22X1 port map( IN1 => addout_49_port, IN2 => n1070, IN3 => 
                           andout_49_port, IN4 => n1059, Q => n697);
   U1476 : AO221X1 port map( IN1 => n51, IN2 => n1092, IN3 => n1081, IN4 => 
                           RAMB(81), IN5 => n697, Q => n698);
   U1477 : OAI21X1 port map( IN1 => n699, IN2 => n698, IN3 => n1136, QN => n701
                           );
   U1478 : OA22X1 port map( IN1 => n1192, IN2 => n1114, IN3 => n1249, IN4 => 
                           n1103, Q => n700);
   U1479 : NAND3X0 port map( IN1 => n701, IN2 => n1123, IN3 => n700, QN => 
                           perm_output(49));
   U1480 : AO22X1 port map( IN1 => eshift_48_port, IN2 => n1026, IN3 => n1015, 
                           IN4 => RAMB(37), Q => n702);
   U1481 : AO221X1 port map( IN1 => n1192, IN2 => n1048, IN3 => n1037, IN4 => 
                           RAMB(48), IN5 => n702, Q => n705);
   U1482 : AO221X1 port map( IN1 => n21, IN2 => n1092, IN3 => n1081, IN4 => 
                           RAMB(80), IN5 => n703, Q => n704);
   U1483 : OAI21X1 port map( IN1 => n705, IN2 => n704, IN3 => n1136, QN => n707
                           );
   U1484 : OA22X1 port map( IN1 => n1191, IN2 => n1114, IN3 => n1248, IN4 => 
                           n1103, Q => n706);
   U1485 : NAND3X0 port map( IN1 => n707, IN2 => n1123, IN3 => n706, QN => 
                           perm_output(48));
   U1486 : AO22X1 port map( IN1 => eshift_47_port, IN2 => n1026, IN3 => n1015, 
                           IN4 => n17, Q => n708);
   U1487 : AO221X1 port map( IN1 => n1191, IN2 => n1048, IN3 => n1037, IN4 => 
                           RAMB(47), IN5 => n708, Q => n711);
   U1488 : AO22X1 port map( IN1 => addout_47_port, IN2 => n1070, IN3 => 
                           andout_47_port, IN4 => n1059, Q => n709);
   U1489 : AO221X1 port map( IN1 => n134, IN2 => n1092, IN3 => n1081, IN4 => 
                           RAMB(79), IN5 => n709, Q => n710);
   U1490 : OAI21X1 port map( IN1 => n711, IN2 => n710, IN3 => n1137, QN => n713
                           );
   U1491 : OA22X1 port map( IN1 => n1190, IN2 => n1114, IN3 => n1247, IN4 => 
                           n1103, Q => n712);
   U1492 : NAND3X0 port map( IN1 => n713, IN2 => n1123, IN3 => n712, QN => 
                           perm_output(47));
   U1493 : AO22X1 port map( IN1 => eshift_46_port, IN2 => n1026, IN3 => n1015, 
                           IN4 => RAMB(35), Q => n714);
   U1494 : AO221X1 port map( IN1 => n1190, IN2 => n1048, IN3 => n1037, IN4 => 
                           RAMB(46), IN5 => n714, Q => n717);
   U1495 : AO22X1 port map( IN1 => addout_46_port, IN2 => n1070, IN3 => 
                           andout_46_port, IN4 => n1059, Q => n715);
   U1496 : AO221X1 port map( IN1 => n85, IN2 => n1092, IN3 => n1081, IN4 => 
                           RAMB(78), IN5 => n715, Q => n716);
   U1497 : OAI21X1 port map( IN1 => n717, IN2 => n716, IN3 => n1137, QN => n719
                           );
   U1498 : OA22X1 port map( IN1 => n1189, IN2 => n1114, IN3 => n1246, IN4 => 
                           n1103, Q => n718);
   U1499 : NAND3X0 port map( IN1 => n719, IN2 => n1123, IN3 => n718, QN => 
                           perm_output(46));
   U1500 : AO22X1 port map( IN1 => eshift_45_port, IN2 => n1026, IN3 => n1015, 
                           IN4 => RAMB(34), Q => n720);
   U1501 : AO221X1 port map( IN1 => n1189, IN2 => n1048, IN3 => n1037, IN4 => 
                           RAMB(45), IN5 => n720, Q => n723);
   U1502 : AO22X1 port map( IN1 => addout_45_port, IN2 => n1070, IN3 => 
                           andout_45_port, IN4 => n1059, Q => n721);
   U1503 : AO221X1 port map( IN1 => n67, IN2 => n1092, IN3 => n1081, IN4 => 
                           RAMB(77), IN5 => n721, Q => n722);
   U1504 : OAI21X1 port map( IN1 => n723, IN2 => n722, IN3 => n1137, QN => n725
                           );
   U1505 : OA22X1 port map( IN1 => n1188, IN2 => n1114, IN3 => n1245, IN4 => 
                           n1103, Q => n724);
   U1506 : NAND3X0 port map( IN1 => n725, IN2 => n1123, IN3 => n724, QN => 
                           perm_output(45));
   U1507 : AO22X1 port map( IN1 => eshift_44_port, IN2 => n1026, IN3 => n1015, 
                           IN4 => RAMB(33), Q => n726);
   U1508 : AO221X1 port map( IN1 => n1188, IN2 => n1048, IN3 => n1037, IN4 => 
                           RAMB(44), IN5 => n726, Q => n729);
   U1509 : AO22X1 port map( IN1 => addout_44_port, IN2 => n1070, IN3 => 
                           andout_44_port, IN4 => n1059, Q => n727);
   U1510 : AO221X1 port map( IN1 => n44, IN2 => n1092, IN3 => n1081, IN4 => 
                           RAMB(76), IN5 => n727, Q => n728);
   U1511 : OAI21X1 port map( IN1 => n729, IN2 => n728, IN3 => n1137, QN => n731
                           );
   U1512 : OA22X1 port map( IN1 => n1187, IN2 => n1114, IN3 => n1244, IN4 => 
                           n1103, Q => n730);
   U1513 : NAND3X0 port map( IN1 => n731, IN2 => n1123, IN3 => n730, QN => 
                           perm_output(44));
   U1514 : AO22X1 port map( IN1 => eshift_43_port, IN2 => n1025, IN3 => n1014, 
                           IN4 => RAMB(32), Q => n732);
   U1515 : AO221X1 port map( IN1 => n1187, IN2 => n1047, IN3 => n1036, IN4 => 
                           RAMB(43), IN5 => n732, Q => n735);
   U1516 : AO22X1 port map( IN1 => addout_43_port, IN2 => n1069, IN3 => 
                           andout_43_port, IN4 => n1058, Q => n733);
   U1517 : AO221X1 port map( IN1 => n40, IN2 => n1091, IN3 => n1080, IN4 => 
                           RAMB(75), IN5 => n733, Q => n734);
   U1518 : OAI21X1 port map( IN1 => n735, IN2 => n734, IN3 => n1137, QN => n737
                           );
   U1519 : OA22X1 port map( IN1 => n1186, IN2 => n1113, IN3 => n1243, IN4 => 
                           n1102, Q => n736);
   U1520 : NAND3X0 port map( IN1 => n737, IN2 => n1122, IN3 => n736, QN => 
                           perm_output(43));
   U1521 : AO22X1 port map( IN1 => eshift_42_port, IN2 => n1025, IN3 => n1014, 
                           IN4 => RAMB(63), Q => n738);
   U1522 : AO221X1 port map( IN1 => n1186, IN2 => n1047, IN3 => n1036, IN4 => 
                           RAMB(42), IN5 => n738, Q => n741);
   U1523 : AO22X1 port map( IN1 => addout_42_port, IN2 => n1069, IN3 => 
                           andout_42_port, IN4 => n1058, Q => n739);
   U1524 : AO221X1 port map( IN1 => n82, IN2 => n1091, IN3 => n1080, IN4 => 
                           RAMB(74), IN5 => n739, Q => n740);
   U1525 : OAI21X1 port map( IN1 => n741, IN2 => n740, IN3 => n1137, QN => n743
                           );
   U1526 : OA22X1 port map( IN1 => n1185, IN2 => n1113, IN3 => n1242, IN4 => 
                           n1102, Q => n742);
   U1527 : NAND3X0 port map( IN1 => n743, IN2 => n1122, IN3 => n742, QN => 
                           perm_output(42));
   U1528 : AO22X1 port map( IN1 => eshift_41_port, IN2 => n1025, IN3 => n1014, 
                           IN4 => RAMB(62), Q => n744);
   U1529 : AO221X1 port map( IN1 => n1185, IN2 => n1047, IN3 => n1036, IN4 => 
                           RAMB(41), IN5 => n744, Q => n747);
   U1530 : AO22X1 port map( IN1 => addout_41_port, IN2 => n1069, IN3 => 
                           andout_41_port, IN4 => n1058, Q => n745);
   U1531 : AO221X1 port map( IN1 => n61, IN2 => n1091, IN3 => n1080, IN4 => 
                           RAMB(73), IN5 => n745, Q => n746);
   U1532 : OAI21X1 port map( IN1 => n747, IN2 => n746, IN3 => n1137, QN => n749
                           );
   U1533 : OA22X1 port map( IN1 => n1184, IN2 => n1113, IN3 => n1241, IN4 => 
                           n1102, Q => n748);
   U1534 : NAND3X0 port map( IN1 => n749, IN2 => n1122, IN3 => n748, QN => 
                           perm_output(41));
   U1535 : AO22X1 port map( IN1 => eshift_40_port, IN2 => n1025, IN3 => n1014, 
                           IN4 => RAMB(61), Q => n750);
   U1536 : AO221X1 port map( IN1 => n1184, IN2 => n1047, IN3 => n1036, IN4 => 
                           RAMB(40), IN5 => n750, Q => n753);
   U1537 : AO22X1 port map( IN1 => addout_40_port, IN2 => n1069, IN3 => 
                           andout_40_port, IN4 => n1058, Q => n751);
   U1538 : AO221X1 port map( IN1 => n74, IN2 => n1091, IN3 => n1080, IN4 => 
                           RAMB(72), IN5 => n751, Q => n752);
   U1539 : OAI21X1 port map( IN1 => n753, IN2 => n752, IN3 => n1137, QN => n755
                           );
   U1540 : OA22X1 port map( IN1 => n1183, IN2 => n1113, IN3 => n1240, IN4 => 
                           n1102, Q => n754);
   U1541 : NAND3X0 port map( IN1 => n755, IN2 => n1122, IN3 => n754, QN => 
                           perm_output(40));
   U1542 : AO22X1 port map( IN1 => eshift_39_port, IN2 => n1025, IN3 => n1014, 
                           IN4 => RAMB(60), Q => n756);
   U1543 : AO221X1 port map( IN1 => n1183, IN2 => n1047, IN3 => n1036, IN4 => 
                           n16, IN5 => n756, Q => n759);
   U1544 : AO22X1 port map( IN1 => addout_39_port, IN2 => n1069, IN3 => 
                           andout_39_port, IN4 => n1058, Q => n757);
   U1545 : AO221X1 port map( IN1 => n64, IN2 => n1091, IN3 => n1080, IN4 => 
                           RAMB(71), IN5 => n757, Q => n758);
   U1546 : OAI21X1 port map( IN1 => n759, IN2 => n758, IN3 => n1137, QN => n761
                           );
   U1547 : OA22X1 port map( IN1 => n1182, IN2 => n1113, IN3 => n1271, IN4 => 
                           n1102, Q => n760);
   U1548 : NAND3X0 port map( IN1 => n761, IN2 => n1122, IN3 => n760, QN => 
                           perm_output(39));
   U1549 : AO22X1 port map( IN1 => eshift_38_port, IN2 => n1025, IN3 => n1014, 
                           IN4 => RAMB(59), Q => n762);
   U1550 : AO221X1 port map( IN1 => n1182, IN2 => n1047, IN3 => n1036, IN4 => 
                           RAMB(38), IN5 => n762, Q => n765);
   U1551 : AO22X1 port map( IN1 => addout_38_port, IN2 => n1069, IN3 => 
                           andout_38_port, IN4 => n1058, Q => n763);
   U1552 : AO221X1 port map( IN1 => n120, IN2 => n1091, IN3 => n1080, IN4 => 
                           RAMB(70), IN5 => n763, Q => n764);
   U1553 : OAI21X1 port map( IN1 => n765, IN2 => n764, IN3 => n1137, QN => n767
                           );
   U1554 : OA22X1 port map( IN1 => n1181, IN2 => n1113, IN3 => n1270, IN4 => 
                           n1102, Q => n766);
   U1555 : NAND3X0 port map( IN1 => n767, IN2 => n1122, IN3 => n766, QN => 
                           perm_output(38));
   U1556 : AO22X1 port map( IN1 => eshift_37_port, IN2 => n1025, IN3 => n1014, 
                           IN4 => RAMB(58), Q => n768);
   U1557 : AO221X1 port map( IN1 => n1181, IN2 => n1047, IN3 => n1036, IN4 => 
                           RAMB(37), IN5 => n768, Q => n771);
   U1558 : AO22X1 port map( IN1 => addout_37_port, IN2 => n1069, IN3 => 
                           andout_37_port, IN4 => n1058, Q => n769);
   U1559 : AO221X1 port map( IN1 => n48, IN2 => n1091, IN3 => n1080, IN4 => 
                           RAMB(69), IN5 => n769, Q => n770);
   U1560 : OAI21X1 port map( IN1 => n771, IN2 => n770, IN3 => n1137, QN => n773
                           );
   U1561 : OA22X1 port map( IN1 => n1180, IN2 => n1113, IN3 => n1269, IN4 => 
                           n1102, Q => n772);
   U1562 : NAND3X0 port map( IN1 => n773, IN2 => n1122, IN3 => n772, QN => 
                           perm_output(37));
   U1563 : AO22X1 port map( IN1 => eshift_36_port, IN2 => n1025, IN3 => n1014, 
                           IN4 => RAMB(57), Q => n774);
   U1564 : AO221X1 port map( IN1 => n1180, IN2 => n1047, IN3 => n1036, IN4 => 
                           n17, IN5 => n774, Q => n777);
   U1565 : AO22X1 port map( IN1 => addout_36_port, IN2 => n1069, IN3 => 
                           andout_36_port, IN4 => n1058, Q => n775);
   U1566 : AO221X1 port map( IN1 => n129, IN2 => n1091, IN3 => n1080, IN4 => 
                           RAMB(68), IN5 => n775, Q => n776);
   U1567 : OAI21X1 port map( IN1 => n777, IN2 => n776, IN3 => n1137, QN => n779
                           );
   U1568 : OA22X1 port map( IN1 => n1179, IN2 => n1113, IN3 => n1268, IN4 => 
                           n1102, Q => n778);
   U1569 : NAND3X0 port map( IN1 => n779, IN2 => n1122, IN3 => n778, QN => 
                           perm_output(36));
   U1570 : AO22X1 port map( IN1 => eshift_35_port, IN2 => n1025, IN3 => n1014, 
                           IN4 => RAMB(56), Q => n780);
   U1571 : AO221X1 port map( IN1 => n1179, IN2 => n1047, IN3 => n1036, IN4 => 
                           RAMB(35), IN5 => n780, Q => n783);
   U1572 : AO22X1 port map( IN1 => addout_35_port, IN2 => n1069, IN3 => 
                           andout_35_port, IN4 => n1058, Q => n781);
   U1573 : AO221X1 port map( IN1 => n99, IN2 => n1091, IN3 => n1080, IN4 => 
                           RAMB(67), IN5 => n781, Q => n782);
   U1574 : OAI21X1 port map( IN1 => n783, IN2 => n782, IN3 => n1138, QN => n785
                           );
   U1575 : OA22X1 port map( IN1 => n1178, IN2 => n1113, IN3 => n1267, IN4 => 
                           n1102, Q => n784);
   U1576 : NAND3X0 port map( IN1 => n785, IN2 => n1122, IN3 => n784, QN => 
                           perm_output(35));
   U1577 : AO22X1 port map( IN1 => eshift_34_port, IN2 => n1025, IN3 => n1014, 
                           IN4 => RAMB(55), Q => n786);
   U1578 : AO221X1 port map( IN1 => n1178, IN2 => n1047, IN3 => n1036, IN4 => 
                           RAMB(34), IN5 => n786, Q => n789);
   U1579 : AO22X1 port map( IN1 => addout_34_port, IN2 => n1069, IN3 => 
                           andout_34_port, IN4 => n1058, Q => n787);
   U1580 : AO221X1 port map( IN1 => n108, IN2 => n1091, IN3 => n1080, IN4 => 
                           RAMB(66), IN5 => n787, Q => n788);
   U1581 : OAI21X1 port map( IN1 => n789, IN2 => n788, IN3 => n1138, QN => n791
                           );
   U1582 : OA22X1 port map( IN1 => n1177, IN2 => n1113, IN3 => n1266, IN4 => 
                           n1102, Q => n790);
   U1583 : NAND3X0 port map( IN1 => n791, IN2 => n1122, IN3 => n790, QN => 
                           perm_output(34));
   U1584 : AO22X1 port map( IN1 => eshift_33_port, IN2 => n1025, IN3 => n1014, 
                           IN4 => RAMB(54), Q => n792);
   U1585 : AO221X1 port map( IN1 => n1177, IN2 => n1047, IN3 => n1036, IN4 => 
                           RAMB(33), IN5 => n792, Q => n795);
   U1586 : AO22X1 port map( IN1 => addout_33_port, IN2 => n1069, IN3 => 
                           andout_33_port, IN4 => n1058, Q => n793);
   U1587 : AO221X1 port map( IN1 => n141, IN2 => n1091, IN3 => n1080, IN4 => 
                           RAMB(65), IN5 => n793, Q => n794);
   U1588 : OAI21X1 port map( IN1 => n795, IN2 => n794, IN3 => n1138, QN => n797
                           );
   U1589 : OA22X1 port map( IN1 => n1176, IN2 => n1113, IN3 => n1265, IN4 => 
                           n1102, Q => n796);
   U1590 : NAND3X0 port map( IN1 => n797, IN2 => n1122, IN3 => n796, QN => 
                           perm_output(33));
   U1591 : AO22X1 port map( IN1 => eshift_32_port, IN2 => n1025, IN3 => n1014, 
                           IN4 => RAMB(53), Q => n798);
   U1592 : AO221X1 port map( IN1 => n1176, IN2 => n1047, IN3 => n1036, IN4 => 
                           RAMB(32), IN5 => n798, Q => n801);
   U1593 : AO22X1 port map( IN1 => addout_32_port, IN2 => n1069, IN3 => 
                           andout_32_port, IN4 => n1058, Q => n799);
   U1594 : AO221X1 port map( IN1 => n83, IN2 => n1091, IN3 => n1080, IN4 => 
                           RAMB(64), IN5 => n799, Q => n800);
   U1595 : OAI21X1 port map( IN1 => n801, IN2 => n800, IN3 => n1138, QN => n803
                           );
   U1596 : OA22X1 port map( IN1 => n1207, IN2 => n1113, IN3 => n1264, IN4 => 
                           n1102, Q => n802);
   U1597 : NAND3X0 port map( IN1 => n803, IN2 => n1122, IN3 => n802, QN => 
                           perm_output(32));
   U1598 : AO22X1 port map( IN1 => eshift_31_port, IN2 => n1024, IN3 => n1013, 
                           IN4 => RAMB(20), Q => n804);
   U1599 : AO221X1 port map( IN1 => n1175, IN2 => n1046, IN3 => n1035, IN4 => 
                           RAMB(31), IN5 => n804, Q => n807);
   U1600 : AO22X1 port map( IN1 => addout_31_port, IN2 => n1068, IN3 => 
                           andout_31_port, IN4 => n1057, Q => n805);
   U1601 : AO221X1 port map( IN1 => n98, IN2 => n1090, IN3 => n1079, IN4 => 
                           RAMB(63), IN5 => n805, Q => n806);
   U1602 : OAI21X1 port map( IN1 => n807, IN2 => n806, IN3 => n1138, QN => n809
                           );
   U1603 : OA22X1 port map( IN1 => n1174, IN2 => n1112, IN3 => n1231, IN4 => 
                           n1101, Q => n808);
   U1604 : NAND3X0 port map( IN1 => n809, IN2 => n1127, IN3 => n808, QN => 
                           perm_output(31));
   U1605 : AO22X1 port map( IN1 => eshift_30_port, IN2 => n1024, IN3 => n1013, 
                           IN4 => RAMB(19), Q => n810);
   U1606 : AO221X1 port map( IN1 => n1174, IN2 => n1046, IN3 => n1035, IN4 => 
                           RAMB(30), IN5 => n810, Q => n813);
   U1607 : AO22X1 port map( IN1 => addout_30_port, IN2 => n1068, IN3 => 
                           andout_30_port, IN4 => n1057, Q => n811);
   U1608 : AO221X1 port map( IN1 => n37, IN2 => n1090, IN3 => n1079, IN4 => 
                           RAMB(62), IN5 => n811, Q => n812);
   U1609 : OAI21X1 port map( IN1 => n813, IN2 => n812, IN3 => n1138, QN => n815
                           );
   U1610 : OA22X1 port map( IN1 => n1173, IN2 => n1112, IN3 => n1230, IN4 => 
                           n1101, Q => n814);
   U1611 : NAND3X0 port map( IN1 => n815, IN2 => n1123, IN3 => n814, QN => 
                           perm_output(30));
   U1612 : AO22X1 port map( IN1 => eshift_29_port, IN2 => n1024, IN3 => n1013, 
                           IN4 => RAMB(18), Q => n816);
   U1613 : AO221X1 port map( IN1 => n1173, IN2 => n1046, IN3 => n1035, IN4 => 
                           RAMB(29), IN5 => n816, Q => n819);
   U1614 : AO22X1 port map( IN1 => addout_29_port, IN2 => n1068, IN3 => 
                           andout_29_port, IN4 => n1057, Q => n817);
   U1615 : AO221X1 port map( IN1 => n126, IN2 => n1090, IN3 => n1079, IN4 => 
                           RAMB(61), IN5 => n817, Q => n818);
   U1616 : OAI21X1 port map( IN1 => n819, IN2 => n818, IN3 => n1138, QN => n821
                           );
   U1617 : OA22X1 port map( IN1 => n1172, IN2 => n1112, IN3 => n1229, IN4 => 
                           n1101, Q => n820);
   U1618 : NAND3X0 port map( IN1 => n821, IN2 => n1122, IN3 => n820, QN => 
                           perm_output(29));
   U1619 : AO22X1 port map( IN1 => eshift_28_port, IN2 => n1024, IN3 => n1013, 
                           IN4 => RAMB(17), Q => n822);
   U1620 : AO221X1 port map( IN1 => n1172, IN2 => n1046, IN3 => n1035, IN4 => 
                           RAMB(28), IN5 => n822, Q => n825);
   U1621 : AO22X1 port map( IN1 => addout_28_port, IN2 => n1068, IN3 => 
                           andout_28_port, IN4 => n1057, Q => n823);
   U1622 : AO221X1 port map( IN1 => n119, IN2 => n1090, IN3 => n1079, IN4 => 
                           RAMB(60), IN5 => n823, Q => n824);
   U1623 : OAI21X1 port map( IN1 => n825, IN2 => n824, IN3 => n1138, QN => n827
                           );
   U1624 : OA22X1 port map( IN1 => n1171, IN2 => n1112, IN3 => n1228, IN4 => 
                           n1101, Q => n826);
   U1625 : NAND3X0 port map( IN1 => n827, IN2 => n1122, IN3 => n826, QN => 
                           perm_output(28));
   U1626 : AO22X1 port map( IN1 => eshift_27_port, IN2 => n1024, IN3 => n1013, 
                           IN4 => RAMB(16), Q => n828);
   U1627 : AO221X1 port map( IN1 => n1171, IN2 => n1046, IN3 => n1035, IN4 => 
                           RAMB(27), IN5 => n828, Q => n831);
   U1628 : AO22X1 port map( IN1 => addout_27_port, IN2 => n1068, IN3 => 
                           andout_27_port, IN4 => n1057, Q => n829);
   U1629 : AO221X1 port map( IN1 => n68, IN2 => n1090, IN3 => n1079, IN4 => 
                           RAMB(59), IN5 => n829, Q => n830);
   U1630 : OAI21X1 port map( IN1 => n831, IN2 => n830, IN3 => n1138, QN => n833
                           );
   U1631 : OA22X1 port map( IN1 => n1170, IN2 => n1112, IN3 => n1227, IN4 => 
                           n1101, Q => n832);
   U1632 : NAND3X0 port map( IN1 => n833, IN2 => n1127, IN3 => n832, QN => 
                           perm_output(27));
   U1633 : AO22X1 port map( IN1 => eshift_26_port, IN2 => n1024, IN3 => n1013, 
                           IN4 => RAMB(15), Q => n834);
   U1634 : AO221X1 port map( IN1 => n1170, IN2 => n1046, IN3 => n1035, IN4 => 
                           RAMB(26), IN5 => n834, Q => n837);
   U1635 : AO22X1 port map( IN1 => addout_26_port, IN2 => n1068, IN3 => 
                           andout_26_port, IN4 => n1057, Q => n835);
   U1636 : AO221X1 port map( IN1 => n205, IN2 => n1090, IN3 => n1079, IN4 => 
                           RAMB(58), IN5 => n835, Q => n836);
   U1637 : OAI21X1 port map( IN1 => n837, IN2 => n836, IN3 => n1138, QN => n839
                           );
   U1638 : OA22X1 port map( IN1 => n1169, IN2 => n1112, IN3 => n1226, IN4 => 
                           n1101, Q => n838);
   U1639 : NAND3X0 port map( IN1 => n839, IN2 => n1121, IN3 => n838, QN => 
                           perm_output(26));
   U1640 : AO22X1 port map( IN1 => eshift_25_port, IN2 => n1024, IN3 => n1013, 
                           IN4 => RAMB(14), Q => n840);
   U1641 : AO221X1 port map( IN1 => n1169, IN2 => n1046, IN3 => n1035, IN4 => 
                           RAMB(25), IN5 => n840, Q => n843);
   U1642 : AO22X1 port map( IN1 => addout_25_port, IN2 => n1068, IN3 => 
                           andout_25_port, IN4 => n1057, Q => n841);
   U1643 : AO221X1 port map( IN1 => n73, IN2 => n1090, IN3 => n1079, IN4 => 
                           RAMB(57), IN5 => n841, Q => n842);
   U1644 : OAI21X1 port map( IN1 => n843, IN2 => n842, IN3 => n1138, QN => n845
                           );
   U1645 : OA22X1 port map( IN1 => n1168, IN2 => n1112, IN3 => n1225, IN4 => 
                           n1101, Q => n844);
   U1646 : NAND3X0 port map( IN1 => n845, IN2 => n1122, IN3 => n844, QN => 
                           perm_output(25));
   U1647 : AO22X1 port map( IN1 => eshift_24_port, IN2 => n1024, IN3 => n1013, 
                           IN4 => RAMB(13), Q => n846);
   U1648 : AO221X1 port map( IN1 => n1168, IN2 => n1046, IN3 => n1035, IN4 => 
                           RAMB(24), IN5 => n846, Q => n849);
   U1649 : AO22X1 port map( IN1 => addout_24_port, IN2 => n1068, IN3 => 
                           andout_24_port, IN4 => n1057, Q => n847);
   U1650 : AO221X1 port map( IN1 => n36, IN2 => n1090, IN3 => n1079, IN4 => 
                           RAMB(56), IN5 => n847, Q => n848);
   U1651 : OAI21X1 port map( IN1 => n849, IN2 => n848, IN3 => n1138, QN => n851
                           );
   U1652 : OA22X1 port map( IN1 => n1167, IN2 => n1112, IN3 => n1224, IN4 => 
                           n1101, Q => n850);
   U1653 : NAND3X0 port map( IN1 => n851, IN2 => n1121, IN3 => n850, QN => 
                           perm_output(24));
   U1654 : AO22X1 port map( IN1 => eshift_23_port, IN2 => n1024, IN3 => n1013, 
                           IN4 => RAMB(12), Q => n852);
   U1655 : AO221X1 port map( IN1 => n1167, IN2 => n1046, IN3 => n1035, IN4 => 
                           RAMB(23), IN5 => n852, Q => n855);
   U1656 : AO22X1 port map( IN1 => addout_23_port, IN2 => n1068, IN3 => 
                           andout_23_port, IN4 => n1057, Q => n853);
   U1657 : AO221X1 port map( IN1 => n43, IN2 => n1090, IN3 => n1079, IN4 => 
                           RAMB(55), IN5 => n853, Q => n854);
   U1658 : OAI21X1 port map( IN1 => n855, IN2 => n854, IN3 => n1139, QN => n857
                           );
   U1659 : OA22X1 port map( IN1 => n1166, IN2 => n1112, IN3 => n1223, IN4 => 
                           n1101, Q => n856);
   U1660 : NAND3X0 port map( IN1 => n857, IN2 => n1123, IN3 => n856, QN => 
                           perm_output(23));
   U1661 : AO22X1 port map( IN1 => eshift_22_port, IN2 => n1024, IN3 => n1013, 
                           IN4 => RAMB(11), Q => n858);
   U1662 : AO221X1 port map( IN1 => n1166, IN2 => n1046, IN3 => n1035, IN4 => 
                           RAMB(22), IN5 => n858, Q => n861);
   U1663 : AO22X1 port map( IN1 => addout_22_port, IN2 => n1068, IN3 => 
                           andout_22_port, IN4 => n1057, Q => n859);
   U1664 : AO221X1 port map( IN1 => n210, IN2 => n1090, IN3 => n1079, IN4 => 
                           RAMB(54), IN5 => n859, Q => n860);
   U1665 : OAI21X1 port map( IN1 => n861, IN2 => n860, IN3 => n1139, QN => n863
                           );
   U1666 : OA22X1 port map( IN1 => n1165, IN2 => n1112, IN3 => n1222, IN4 => 
                           n1101, Q => n862);
   U1667 : AO22X1 port map( IN1 => eshift_21_port, IN2 => n1024, IN3 => n1013, 
                           IN4 => RAMB(10), Q => n864);
   U1668 : AO221X1 port map( IN1 => n1165, IN2 => n1046, IN3 => n1035, IN4 => 
                           RAMB(21), IN5 => n864, Q => n867);
   U1669 : AO22X1 port map( IN1 => addout_21_port, IN2 => n1068, IN3 => 
                           andout_21_port, IN4 => n1057, Q => n865);
   U1670 : AO221X1 port map( IN1 => n201, IN2 => n1090, IN3 => n1079, IN4 => 
                           RAMB(53), IN5 => n865, Q => n866);
   U1671 : OAI21X1 port map( IN1 => n867, IN2 => n866, IN3 => n1139, QN => n869
                           );
   U1672 : OA22X1 port map( IN1 => n1164, IN2 => n1112, IN3 => n1221, IN4 => 
                           n1101, Q => n868);
   U1673 : NAND3X0 port map( IN1 => n869, IN2 => n1127, IN3 => n868, QN => 
                           perm_output(21));
   U1674 : AO22X1 port map( IN1 => eshift_20_port, IN2 => n1024, IN3 => n1013, 
                           IN4 => RAMB(9), Q => n870);
   U1675 : AO221X1 port map( IN1 => n1164, IN2 => n1046, IN3 => n1035, IN4 => 
                           RAMB(20), IN5 => n870, Q => n873);
   U1676 : AO22X1 port map( IN1 => addout_20_port, IN2 => n1068, IN3 => 
                           andout_20_port, IN4 => n1057, Q => n871);
   U1677 : AO221X1 port map( IN1 => n132, IN2 => n1090, IN3 => n1079, IN4 => 
                           RAMB(52), IN5 => n871, Q => n872);
   U1678 : OAI21X1 port map( IN1 => n873, IN2 => n872, IN3 => n1139, QN => n875
                           );
   U1679 : OA22X1 port map( IN1 => n1163, IN2 => n1112, IN3 => n1220, IN4 => 
                           n1101, Q => n874);
   U1680 : NAND3X0 port map( IN1 => n875, IN2 => n1128, IN3 => n874, QN => 
                           perm_output(20));
   U1681 : AO22X1 port map( IN1 => eshift_19_port, IN2 => n1023, IN3 => n1012, 
                           IN4 => RAMB(8), Q => n876);
   U1682 : AO221X1 port map( IN1 => n1163, IN2 => n1045, IN3 => n1034, IN4 => 
                           RAMB(19), IN5 => n876, Q => n879);
   U1683 : AO22X1 port map( IN1 => addout_19_port, IN2 => n1067, IN3 => 
                           andout_19_port, IN4 => n1056, Q => n877);
   U1684 : AO221X1 port map( IN1 => n72, IN2 => n1089, IN3 => n1078, IN4 => 
                           RAMB(51), IN5 => n877, Q => n878);
   U1685 : OAI21X1 port map( IN1 => n879, IN2 => n878, IN3 => n1139, QN => n881
                           );
   U1686 : OA22X1 port map( IN1 => n1162, IN2 => n1111, IN3 => n1219, IN4 => 
                           n1100, Q => n880);
   U1687 : NAND3X0 port map( IN1 => n881, IN2 => n1121, IN3 => n880, QN => 
                           perm_output(19));
   U1688 : AO22X1 port map( IN1 => eshift_18_port, IN2 => n1023, IN3 => n1012, 
                           IN4 => RAMB(7), Q => n882);
   U1689 : AO221X1 port map( IN1 => n1162, IN2 => n1045, IN3 => n1034, IN4 => 
                           RAMB(18), IN5 => n882, Q => n885);
   U1690 : AO22X1 port map( IN1 => addout_18_port, IN2 => n1067, IN3 => 
                           andout_18_port, IN4 => n1056, Q => n883);
   U1691 : AO221X1 port map( IN1 => n55, IN2 => n1089, IN3 => n1078, IN4 => 
                           RAMB(50), IN5 => n883, Q => n884);
   U1692 : OAI21X1 port map( IN1 => n885, IN2 => n884, IN3 => n1139, QN => n887
                           );
   U1693 : OA22X1 port map( IN1 => n1161, IN2 => n1111, IN3 => n1218, IN4 => 
                           n1100, Q => n886);
   U1694 : NAND3X0 port map( IN1 => n887, IN2 => n1121, IN3 => n886, QN => 
                           perm_output(18));
   U1695 : AO22X1 port map( IN1 => eshift_17_port, IN2 => n1023, IN3 => n1012, 
                           IN4 => RAMB(6), Q => n888);
   U1696 : AO221X1 port map( IN1 => n1161, IN2 => n1045, IN3 => n1034, IN4 => 
                           RAMB(17), IN5 => n888, Q => n891);
   U1697 : AO22X1 port map( IN1 => addout_17_port, IN2 => n1067, IN3 => 
                           andout_17_port, IN4 => n1056, Q => n889);
   U1698 : AO221X1 port map( IN1 => n122, IN2 => n1089, IN3 => n1078, IN4 => 
                           RAMB(49), IN5 => n889, Q => n890);
   U1699 : OAI21X1 port map( IN1 => n891, IN2 => n890, IN3 => n1139, QN => n893
                           );
   U1700 : OA22X1 port map( IN1 => n1160, IN2 => n1111, IN3 => n1217, IN4 => 
                           n1100, Q => n892);
   U1701 : NAND3X0 port map( IN1 => n893, IN2 => n1121, IN3 => n892, QN => 
                           perm_output(17));
   U1702 : AO22X1 port map( IN1 => eshift_16_port, IN2 => n1023, IN3 => n1012, 
                           IN4 => RAMB(5), Q => n894);
   U1703 : AO221X1 port map( IN1 => n1160, IN2 => n1045, IN3 => n1034, IN4 => 
                           RAMB(16), IN5 => n894, Q => n897);
   U1704 : AO22X1 port map( IN1 => addout_16_port, IN2 => n1067, IN3 => 
                           andout_16_port, IN4 => n1056, Q => n895);
   U1705 : AO221X1 port map( IN1 => n117, IN2 => n1089, IN3 => n1078, IN4 => 
                           RAMB(48), IN5 => n895, Q => n896);
   U1706 : OAI21X1 port map( IN1 => n897, IN2 => n896, IN3 => n1139, QN => n899
                           );
   U1707 : OA22X1 port map( IN1 => n1159, IN2 => n1111, IN3 => n1216, IN4 => 
                           n1100, Q => n898);
   U1708 : NAND3X0 port map( IN1 => n899, IN2 => n1121, IN3 => n898, QN => 
                           perm_output(16));
   U1709 : AO22X1 port map( IN1 => eshift_15_port, IN2 => n1023, IN3 => n1012, 
                           IN4 => RAMB(4), Q => n900);
   U1710 : AO221X1 port map( IN1 => n1159, IN2 => n1045, IN3 => n1034, IN4 => 
                           RAMB(15), IN5 => n900, Q => n903);
   U1711 : AO22X1 port map( IN1 => addout_15_port, IN2 => n1067, IN3 => 
                           andout_15_port, IN4 => n1056, Q => n901);
   U1712 : AO221X1 port map( IN1 => n101, IN2 => n1089, IN3 => n1078, IN4 => 
                           RAMB(47), IN5 => n901, Q => n902);
   U1713 : OAI21X1 port map( IN1 => n903, IN2 => n902, IN3 => n1139, QN => n905
                           );
   U1714 : OA22X1 port map( IN1 => n1158, IN2 => n1111, IN3 => n1215, IN4 => 
                           n1100, Q => n904);
   U1715 : NAND3X0 port map( IN1 => n905, IN2 => n1121, IN3 => n904, QN => 
                           perm_output(15));
   U1716 : AO22X1 port map( IN1 => eshift_14_port, IN2 => n1023, IN3 => n1012, 
                           IN4 => RAMB(3), Q => n906);
   U1717 : AO221X1 port map( IN1 => n1158, IN2 => n1045, IN3 => n1034, IN4 => 
                           RAMB(14), IN5 => n906, Q => n909);
   U1718 : AO22X1 port map( IN1 => addout_14_port, IN2 => n1067, IN3 => 
                           andout_14_port, IN4 => n1056, Q => n907);
   U1719 : AO221X1 port map( IN1 => n125, IN2 => n1089, IN3 => n1078, IN4 => 
                           RAMB(46), IN5 => n907, Q => n908);
   U1720 : OAI21X1 port map( IN1 => n909, IN2 => n908, IN3 => n1139, QN => n911
                           );
   U1721 : OA22X1 port map( IN1 => n1157, IN2 => n1111, IN3 => n1214, IN4 => 
                           n1100, Q => n910);
   U1722 : NAND3X0 port map( IN1 => n911, IN2 => n1121, IN3 => n910, QN => 
                           perm_output(14));
   U1723 : AO22X1 port map( IN1 => eshift_13_port, IN2 => n1023, IN3 => n1012, 
                           IN4 => RAMB(2), Q => n912);
   U1724 : AO221X1 port map( IN1 => n1157, IN2 => n1045, IN3 => n1034, IN4 => 
                           RAMB(13), IN5 => n912, Q => n915);
   U1725 : AO22X1 port map( IN1 => addout_13_port, IN2 => n1067, IN3 => 
                           andout_13_port, IN4 => n1056, Q => n913);
   U1726 : AO221X1 port map( IN1 => n127, IN2 => n1089, IN3 => n1078, IN4 => 
                           RAMB(45), IN5 => n913, Q => n914);
   U1727 : OAI21X1 port map( IN1 => n915, IN2 => n914, IN3 => n1139, QN => n917
                           );
   U1728 : OA22X1 port map( IN1 => n1156, IN2 => n1111, IN3 => n1213, IN4 => 
                           n1100, Q => n916);
   U1729 : NAND3X0 port map( IN1 => n917, IN2 => n1121, IN3 => n916, QN => 
                           perm_output(13));
   U1730 : AO22X1 port map( IN1 => eshift_12_port, IN2 => n1023, IN3 => n1012, 
                           IN4 => RAMB(1), Q => n918);
   U1731 : AO221X1 port map( IN1 => n1156, IN2 => n1045, IN3 => n1034, IN4 => 
                           RAMB(12), IN5 => n918, Q => n921);
   U1732 : AO22X1 port map( IN1 => addout_12_port, IN2 => n1067, IN3 => 
                           andout_12_port, IN4 => n1056, Q => n919);
   U1733 : AO221X1 port map( IN1 => n75, IN2 => n1089, IN3 => n1078, IN4 => 
                           RAMB(44), IN5 => n919, Q => n920);
   U1734 : OAI21X1 port map( IN1 => n921, IN2 => n920, IN3 => n1139, QN => n923
                           );
   U1735 : OA22X1 port map( IN1 => n1155, IN2 => n1111, IN3 => n1212, IN4 => 
                           n1100, Q => n922);
   U1736 : NAND3X0 port map( IN1 => n923, IN2 => n1121, IN3 => n922, QN => 
                           perm_output(12));
   U1737 : AO22X1 port map( IN1 => eshift_11_port, IN2 => n1023, IN3 => n1012, 
                           IN4 => RAMB(0), Q => n924);
   U1738 : AO221X1 port map( IN1 => n1155, IN2 => n1045, IN3 => n1034, IN4 => 
                           RAMB(11), IN5 => n924, Q => n927);
   U1739 : AO22X1 port map( IN1 => addout_11_port, IN2 => n1067, IN3 => 
                           andout_11_port, IN4 => n1056, Q => n925);
   U1740 : AO221X1 port map( IN1 => n97, IN2 => n1089, IN3 => n1078, IN4 => 
                           RAMB(43), IN5 => n925, Q => n926);
   U1741 : OAI21X1 port map( IN1 => n927, IN2 => n926, IN3 => n1140, QN => n929
                           );
   U1742 : OA22X1 port map( IN1 => n1154, IN2 => n1111, IN3 => n1211, IN4 => 
                           n1100, Q => n928);
   U1743 : NAND3X0 port map( IN1 => n929, IN2 => n1121, IN3 => n928, QN => 
                           perm_output(11));
   U1744 : AO22X1 port map( IN1 => eshift_10_port, IN2 => n1023, IN3 => n1012, 
                           IN4 => RAMB(31), Q => n930);
   U1745 : AO221X1 port map( IN1 => n1154, IN2 => n1045, IN3 => n1034, IN4 => 
                           RAMB(10), IN5 => n930, Q => n933);
   U1746 : AO22X1 port map( IN1 => n1067, IN2 => addout_10_port, IN3 => 
                           andout_10_port, IN4 => n1056, Q => n931);
   U1747 : AO221X1 port map( IN1 => n93, IN2 => n1089, IN3 => n1078, IN4 => 
                           RAMB(42), IN5 => n931, Q => n932);
   U1748 : OAI21X1 port map( IN1 => n933, IN2 => n932, IN3 => n1140, QN => n935
                           );
   U1749 : OA22X1 port map( IN1 => n1153, IN2 => n1111, IN3 => n1210, IN4 => 
                           n1100, Q => n934);
   U1750 : NAND3X0 port map( IN1 => n935, IN2 => n1121, IN3 => n934, QN => 
                           perm_output(10));
   U1751 : AO22X1 port map( IN1 => eshift_9_port, IN2 => n1023, IN3 => n1012, 
                           IN4 => RAMB(30), Q => n936);
   U1752 : AO221X1 port map( IN1 => n1153, IN2 => n1045, IN3 => n1034, IN4 => 
                           RAMB(9), IN5 => n936, Q => n939);
   U1753 : AO22X1 port map( IN1 => addout_9_port, IN2 => n1067, IN3 => 
                           andout_9_port, IN4 => n1056, Q => n937);
   U1754 : AO221X1 port map( IN1 => n92, IN2 => n1089, IN3 => n1078, IN4 => 
                           RAMB(41), IN5 => n937, Q => n938);
   U1755 : OAI21X1 port map( IN1 => n939, IN2 => n938, IN3 => n1140, QN => n941
                           );
   U1756 : OA22X1 port map( IN1 => n1152, IN2 => n1111, IN3 => n1209, IN4 => 
                           n1100, Q => n940);
   U1757 : NAND3X0 port map( IN1 => n941, IN2 => n1121, IN3 => n940, QN => 
                           perm_output(9));
   U1758 : AO22X1 port map( IN1 => eshift_8_port, IN2 => n1023, IN3 => n1012, 
                           IN4 => RAMB(29), Q => n942);
   U1759 : AO221X1 port map( IN1 => n1152, IN2 => n1045, IN3 => n1034, IN4 => 
                           RAMB(8), IN5 => n942, Q => n945);
   U1760 : AO22X1 port map( IN1 => addout_8_port, IN2 => n1067, IN3 => 
                           andout_8_port, IN4 => n1056, Q => n943);
   U1761 : AO221X1 port map( IN1 => n102, IN2 => n1089, IN3 => n1078, IN4 => 
                           RAMB(40), IN5 => n943, Q => n944);
   U1762 : OAI21X1 port map( IN1 => n945, IN2 => n944, IN3 => n1140, QN => n947
                           );
   U1763 : OA22X1 port map( IN1 => n1151, IN2 => n1111, IN3 => n1208, IN4 => 
                           n1100, Q => n946);
   U1764 : NAND3X0 port map( IN1 => n947, IN2 => n1121, IN3 => n946, QN => 
                           perm_output(8));
   U1765 : AO22X1 port map( IN1 => eshift_7_port, IN2 => n1022, IN3 => n1011, 
                           IN4 => RAMB(28), Q => n948);
   U1766 : AO221X1 port map( IN1 => n1151, IN2 => n1044, IN3 => n1033, IN4 => 
                           RAMB(7), IN5 => n948, Q => n951);
   U1767 : AO22X1 port map( IN1 => addout_7_port, IN2 => n1066, IN3 => 
                           andout_7_port, IN4 => n1055, Q => n949);
   U1768 : AO221X1 port map( IN1 => n111, IN2 => n1088, IN3 => n1077, IN4 => 
                           n16, IN5 => n949, Q => n950);
   U1769 : OAI21X1 port map( IN1 => n951, IN2 => n950, IN3 => n1140, QN => n953
                           );
   U1770 : OA22X1 port map( IN1 => n1150, IN2 => n1110, IN3 => n1239, IN4 => 
                           n1099, Q => n952);
   U1771 : AO22X1 port map( IN1 => eshift_6_port, IN2 => n1022, IN3 => n1011, 
                           IN4 => RAMB(27), Q => n954);
   U1772 : AO221X1 port map( IN1 => n1150, IN2 => n1044, IN3 => n1033, IN4 => 
                           RAMB(6), IN5 => n954, Q => n957);
   U1773 : AO22X1 port map( IN1 => addout_6_port, IN2 => n1066, IN3 => 
                           andout_6_port, IN4 => n1055, Q => n955);
   U1774 : AO221X1 port map( IN1 => n135, IN2 => n1088, IN3 => n1077, IN4 => 
                           RAMB(38), IN5 => n955, Q => n956);
   U1775 : OAI21X1 port map( IN1 => n957, IN2 => n956, IN3 => n1140, QN => n959
                           );
   U1776 : OA22X1 port map( IN1 => n1149, IN2 => n1110, IN3 => n1238, IN4 => 
                           n1099, Q => n958);
   U1777 : NAND3X0 port map( IN1 => n959, IN2 => n1128, IN3 => n958, QN => 
                           perm_output(6));
   U1778 : AO22X1 port map( IN1 => eshift_5_port, IN2 => n1022, IN3 => n1011, 
                           IN4 => RAMB(26), Q => n960);
   U1779 : AO221X1 port map( IN1 => n1149, IN2 => n1044, IN3 => n1033, IN4 => 
                           RAMB(5), IN5 => n960, Q => n963);
   U1780 : AO22X1 port map( IN1 => addout_5_port, IN2 => n1066, IN3 => 
                           andout_5_port, IN4 => n1055, Q => n961);
   U1781 : AO221X1 port map( IN1 => n60, IN2 => n1088, IN3 => n1077, IN4 => 
                           RAMB(37), IN5 => n961, Q => n962);
   U1782 : OAI21X1 port map( IN1 => n963, IN2 => n962, IN3 => n1140, QN => n965
                           );
   U1783 : OA22X1 port map( IN1 => n1148, IN2 => n1110, IN3 => n1237, IN4 => 
                           n1099, Q => n964);
   U1784 : NAND3X0 port map( IN1 => n965, IN2 => n1122, IN3 => n964, QN => 
                           perm_output(5));
   U1785 : AO22X1 port map( IN1 => eshift_4_port, IN2 => n1022, IN3 => n1011, 
                           IN4 => RAMB(25), Q => n966);
   U1786 : AO221X1 port map( IN1 => n1148, IN2 => n1044, IN3 => n1033, IN4 => 
                           RAMB(4), IN5 => n966, Q => n969);
   U1787 : AO22X1 port map( IN1 => addout_4_port, IN2 => n1066, IN3 => 
                           andout_4_port, IN4 => n1055, Q => n967);
   U1788 : AO221X1 port map( IN1 => n89, IN2 => n1088, IN3 => n1077, IN4 => n17
                           , IN5 => n967, Q => n968);
   U1789 : OAI21X1 port map( IN1 => n969, IN2 => n968, IN3 => n1140, QN => n971
                           );
   U1790 : OA22X1 port map( IN1 => n1147, IN2 => n1110, IN3 => n1236, IN4 => 
                           n1099, Q => n970);
   U1791 : NAND3X0 port map( IN1 => n971, IN2 => n1123, IN3 => n970, QN => 
                           perm_output(4));
   U1792 : AO22X1 port map( IN1 => eshift_3_port, IN2 => n1022, IN3 => n1011, 
                           IN4 => RAMB(24), Q => n972);
   U1793 : AO221X1 port map( IN1 => n1147, IN2 => n1044, IN3 => n1033, IN4 => 
                           RAMB(3), IN5 => n972, Q => n975);
   U1794 : AO22X1 port map( IN1 => addout_3_port, IN2 => n1066, IN3 => 
                           andout_3_port, IN4 => n1055, Q => n973);
   U1795 : AO221X1 port map( IN1 => n59, IN2 => n1088, IN3 => n1077, IN4 => 
                           RAMB(35), IN5 => n973, Q => n974);
   U1796 : OAI21X1 port map( IN1 => n975, IN2 => n974, IN3 => n1140, QN => n977
                           );
   U1797 : OA22X1 port map( IN1 => n1146, IN2 => n1110, IN3 => n1235, IN4 => 
                           n1099, Q => n976);
   U1798 : NAND3X0 port map( IN1 => n977, IN2 => n1127, IN3 => n976, QN => 
                           perm_output(3));
   U1799 : AO22X1 port map( IN1 => eshift_2_port, IN2 => n1022, IN3 => n1011, 
                           IN4 => RAMB(23), Q => n978);
   U1800 : AO221X1 port map( IN1 => n1146, IN2 => n1044, IN3 => n1033, IN4 => 
                           RAMB(2), IN5 => n978, Q => n981);
   U1801 : AO22X1 port map( IN1 => addout_2_port, IN2 => n1066, IN3 => 
                           andout_2_port, IN4 => n1055, Q => n979);
   U1802 : AO221X1 port map( IN1 => n208, IN2 => n1088, IN3 => n1077, IN4 => 
                           RAMB(34), IN5 => n979, Q => n980);
   U1803 : OAI21X1 port map( IN1 => n981, IN2 => n980, IN3 => n1140, QN => n983
                           );
   U1804 : OA22X1 port map( IN1 => n1145, IN2 => n1110, IN3 => n1234, IN4 => 
                           n1099, Q => n982);
   U1805 : NAND3X0 port map( IN1 => n983, IN2 => n1128, IN3 => n982, QN => 
                           perm_output(2));
   U1806 : AO22X1 port map( IN1 => eshift_1_port, IN2 => n1022, IN3 => n1011, 
                           IN4 => RAMB(22), Q => n984);
   U1807 : AO221X1 port map( IN1 => n1145, IN2 => n1044, IN3 => n1033, IN4 => 
                           RAMB(1), IN5 => n984, Q => n987);
   U1808 : AO22X1 port map( IN1 => addout_1_port, IN2 => n1066, IN3 => 
                           andout_1_port, IN4 => n1055, Q => n985);
   U1809 : AO221X1 port map( IN1 => n130, IN2 => n1088, IN3 => n1077, IN4 => 
                           RAMB(33), IN5 => n985, Q => n986);
   U1810 : OAI21X1 port map( IN1 => n987, IN2 => n986, IN3 => n1140, QN => n989
                           );
   U1811 : OA22X1 port map( IN1 => n1144, IN2 => n1110, IN3 => n1233, IN4 => 
                           n1099, Q => n988);
   U1812 : NAND3X0 port map( IN1 => n989, IN2 => n1121, IN3 => n988, QN => 
                           perm_output(1));
   U1813 : AO22X1 port map( IN1 => eshift_0_port, IN2 => n1022, IN3 => n1011, 
                           IN4 => RAMB(21), Q => n992);
   U1814 : AO221X1 port map( IN1 => n1144, IN2 => n1044, IN3 => n1033, IN4 => 
                           RAMB(0), IN5 => n992, Q => n1001);
   U1815 : AO22X1 port map( IN1 => addout_0_port, IN2 => n1066, IN3 => 
                           andout_0_port, IN4 => n1055, Q => n997);
   U1816 : AO221X1 port map( IN1 => n84, IN2 => n1088, IN3 => n1077, IN4 => 
                           RAMB(32), IN5 => n997, Q => n1000);
   U1817 : OAI21X1 port map( IN1 => n1001, IN2 => n1000, IN3 => n1140, QN => 
                           n1006);
   U1818 : OA22X1 port map( IN1 => n1175, IN2 => n1110, IN3 => n1232, IN4 => 
                           n1099, Q => n1004);
   U1819 : NAND3X0 port map( IN1 => n1006, IN2 => n1121, IN3 => n1004, QN => 
                           perm_output(0));
   U1820 : NAND2X1 port map( IN1 => instruction_11_port, IN2 => n231, QN => 
                           n1005);
   U1821 : NAND2X1 port map( IN1 => instruction_11_port, IN2 => n1009, QN => 
                           n1003);
   U1822 : NAND2X1 port map( IN1 => instruction_11_port, IN2 => 
                           instruction_8_port, QN => n1002);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_LWC_1.all;

entity DUAL_PORT_RAM_32_BIT_ADDRESS_LEN128_ADDR_ENTRIES16_ADD_ENT_BITS4_1 is

   port( RAMADDR1, RAMADDR2 : in std_logic_vector (3 downto 0);  RAMDIN1 : in 
         std_logic_vector (127 downto 0);  RAMDOUT1, RAMDOUT2 : out 
         std_logic_vector (127 downto 0);  RAMWRITE1, clk : in std_logic);

end DUAL_PORT_RAM_32_BIT_ADDRESS_LEN128_ADDR_ENTRIES16_ADD_ENT_BITS4_1;

architecture SYN_Behavioral of 
   DUAL_PORT_RAM_32_BIT_ADDRESS_LEN128_ADDR_ENTRIES16_ADD_ENT_BITS4_1 is

   component NOR2X0
      port( IN1, IN2 : in std_logic;  QN : out std_logic);
   end component;
   
   component NAND2X0
      port( IN1, IN2 : in std_logic;  QN : out std_logic);
   end component;
   
   component INVX0
      port( INP : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2X1
      port( IN1, IN2 : in std_logic;  Q : out std_logic);
   end component;
   
   component AND2X2
      port( IN1, IN2 : in std_logic;  Q : out std_logic);
   end component;
   
   component OR4X1
      port( IN1, IN2, IN3, IN4 : in std_logic;  Q : out std_logic);
   end component;
   
   component AO221X1
      port( IN1, IN2, IN3, IN4, IN5 : in std_logic;  Q : out std_logic);
   end component;
   
   component AO22X1
      port( IN1, IN2, IN3, IN4 : in std_logic;  Q : out std_logic);
   end component;
   
   component NBUFFX2
      port( INP : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI221X1
      port( IN1, IN2, IN3, IN4, IN5 : in std_logic;  QN : out std_logic);
   end component;
   
   component NAND4X0
      port( IN1, IN2, IN3, IN4 : in std_logic;  QN : out std_logic);
   end component;
   
   component DELLN1X2
      port( INP : in std_logic;  Z : out std_logic);
   end component;
   
   component AO22X2
      port( IN1, IN2, IN3, IN4 : in std_logic;  Q : out std_logic);
   end component;
   
   component AND2X4
      port( IN1, IN2 : in std_logic;  Q : out std_logic);
   end component;
   
   component IBUFFX16
      port( INP : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221X2
      port( IN1, IN2, IN3, IN4, IN5 : in std_logic;  QN : out std_logic);
   end component;
   
   component OR4X2
      port( IN1, IN2, IN3, IN4 : in std_logic;  Q : out std_logic);
   end component;
   
   component DELLN2X2
      port( INP : in std_logic;  Z : out std_logic);
   end component;
   
   component AO221X2
      port( IN1, IN2, IN3, IN4, IN5 : in std_logic;  Q : out std_logic);
   end component;
   
   component NBUFFX4
      port( INP : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFX1
      port( D, CLK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal RAM_0_127_port, RAM_0_126_port, RAM_0_125_port, RAM_0_124_port, 
      RAM_0_123_port, RAM_0_122_port, RAM_0_121_port, RAM_0_120_port, 
      RAM_0_119_port, RAM_0_118_port, RAM_0_117_port, RAM_0_116_port, 
      RAM_0_115_port, RAM_0_114_port, RAM_0_113_port, RAM_0_112_port, 
      RAM_0_111_port, RAM_0_110_port, RAM_0_109_port, RAM_0_108_port, 
      RAM_0_107_port, RAM_0_106_port, RAM_0_105_port, RAM_0_104_port, 
      RAM_0_103_port, RAM_0_102_port, RAM_0_101_port, RAM_0_100_port, 
      RAM_0_99_port, RAM_0_98_port, RAM_0_97_port, RAM_0_96_port, RAM_0_95_port
      , RAM_0_94_port, RAM_0_93_port, RAM_0_92_port, RAM_0_91_port, 
      RAM_0_90_port, RAM_0_89_port, RAM_0_88_port, RAM_0_87_port, RAM_0_86_port
      , RAM_0_85_port, RAM_0_84_port, RAM_0_83_port, RAM_0_82_port, 
      RAM_0_81_port, RAM_0_80_port, RAM_0_79_port, RAM_0_78_port, RAM_0_77_port
      , RAM_0_76_port, RAM_0_75_port, RAM_0_74_port, RAM_0_73_port, 
      RAM_0_72_port, RAM_0_71_port, RAM_0_70_port, RAM_0_69_port, RAM_0_68_port
      , RAM_0_67_port, RAM_0_66_port, RAM_0_65_port, RAM_0_64_port, 
      RAM_0_63_port, RAM_0_62_port, RAM_0_61_port, RAM_0_60_port, RAM_0_59_port
      , RAM_0_58_port, RAM_0_57_port, RAM_0_56_port, RAM_0_55_port, 
      RAM_0_54_port, RAM_0_53_port, RAM_0_52_port, RAM_0_51_port, RAM_0_50_port
      , RAM_0_49_port, RAM_0_48_port, RAM_0_47_port, RAM_0_46_port, 
      RAM_0_45_port, RAM_0_44_port, RAM_0_43_port, RAM_0_42_port, RAM_0_41_port
      , RAM_0_40_port, RAM_0_39_port, RAM_0_38_port, RAM_0_37_port, 
      RAM_0_36_port, RAM_0_35_port, RAM_0_34_port, RAM_0_33_port, RAM_0_32_port
      , RAM_0_31_port, RAM_0_30_port, RAM_0_29_port, RAM_0_28_port, 
      RAM_0_27_port, RAM_0_26_port, RAM_0_25_port, RAM_0_24_port, RAM_0_23_port
      , RAM_0_22_port, RAM_0_21_port, RAM_0_20_port, RAM_0_19_port, 
      RAM_0_18_port, RAM_0_17_port, RAM_0_16_port, RAM_0_15_port, RAM_0_14_port
      , RAM_0_13_port, RAM_0_12_port, RAM_0_11_port, RAM_0_10_port, 
      RAM_0_9_port, RAM_0_8_port, RAM_0_7_port, RAM_0_6_port, RAM_0_5_port, 
      RAM_0_4_port, RAM_0_3_port, RAM_0_2_port, RAM_0_1_port, RAM_0_0_port, 
      RAM_1_127_port, RAM_1_126_port, RAM_1_125_port, RAM_1_124_port, 
      RAM_1_123_port, RAM_1_122_port, RAM_1_121_port, RAM_1_120_port, 
      RAM_1_119_port, RAM_1_118_port, RAM_1_117_port, RAM_1_116_port, 
      RAM_1_115_port, RAM_1_114_port, RAM_1_113_port, RAM_1_112_port, 
      RAM_1_111_port, RAM_1_110_port, RAM_1_109_port, RAM_1_108_port, 
      RAM_1_107_port, RAM_1_106_port, RAM_1_105_port, RAM_1_104_port, 
      RAM_1_103_port, RAM_1_102_port, RAM_1_101_port, RAM_1_100_port, 
      RAM_1_99_port, RAM_1_98_port, RAM_1_97_port, RAM_1_96_port, RAM_1_95_port
      , RAM_1_94_port, RAM_1_93_port, RAM_1_92_port, RAM_1_91_port, 
      RAM_1_90_port, RAM_1_89_port, RAM_1_88_port, RAM_1_87_port, RAM_1_86_port
      , RAM_1_85_port, RAM_1_84_port, RAM_1_83_port, RAM_1_82_port, 
      RAM_1_81_port, RAM_1_80_port, RAM_1_79_port, RAM_1_78_port, RAM_1_77_port
      , RAM_1_76_port, RAM_1_75_port, RAM_1_74_port, RAM_1_73_port, 
      RAM_1_72_port, RAM_1_71_port, RAM_1_70_port, RAM_1_69_port, RAM_1_68_port
      , RAM_1_67_port, RAM_1_66_port, RAM_1_65_port, RAM_1_64_port, 
      RAM_1_63_port, RAM_1_62_port, RAM_1_61_port, RAM_1_60_port, RAM_1_59_port
      , RAM_1_58_port, RAM_1_57_port, RAM_1_56_port, RAM_1_55_port, 
      RAM_1_54_port, RAM_1_53_port, RAM_1_52_port, RAM_1_51_port, RAM_1_50_port
      , RAM_1_49_port, RAM_1_48_port, RAM_1_47_port, RAM_1_46_port, 
      RAM_1_45_port, RAM_1_44_port, RAM_1_43_port, RAM_1_42_port, RAM_1_41_port
      , RAM_1_40_port, RAM_1_39_port, RAM_1_38_port, RAM_1_37_port, 
      RAM_1_36_port, RAM_1_35_port, RAM_1_34_port, RAM_1_33_port, RAM_1_32_port
      , RAM_1_31_port, RAM_1_30_port, RAM_1_29_port, RAM_1_28_port, 
      RAM_1_27_port, RAM_1_26_port, RAM_1_25_port, RAM_1_24_port, RAM_1_23_port
      , RAM_1_22_port, RAM_1_21_port, RAM_1_20_port, RAM_1_19_port, 
      RAM_1_18_port, RAM_1_17_port, RAM_1_16_port, RAM_1_15_port, RAM_1_14_port
      , RAM_1_13_port, RAM_1_12_port, RAM_1_11_port, RAM_1_10_port, 
      RAM_1_9_port, RAM_1_8_port, RAM_1_7_port, RAM_1_6_port, RAM_1_5_port, 
      RAM_1_4_port, RAM_1_3_port, RAM_1_2_port, RAM_1_1_port, RAM_1_0_port, 
      RAM_2_127_port, RAM_2_126_port, RAM_2_125_port, RAM_2_124_port, 
      RAM_2_123_port, RAM_2_122_port, RAM_2_121_port, RAM_2_120_port, 
      RAM_2_119_port, RAM_2_118_port, RAM_2_117_port, RAM_2_116_port, 
      RAM_2_115_port, RAM_2_114_port, RAM_2_113_port, RAM_2_112_port, 
      RAM_2_111_port, RAM_2_110_port, RAM_2_109_port, RAM_2_108_port, 
      RAM_2_107_port, RAM_2_106_port, RAM_2_105_port, RAM_2_104_port, 
      RAM_2_103_port, RAM_2_102_port, RAM_2_101_port, RAM_2_100_port, 
      RAM_2_99_port, RAM_2_98_port, RAM_2_97_port, RAM_2_96_port, RAM_2_95_port
      , RAM_2_94_port, RAM_2_93_port, RAM_2_92_port, RAM_2_91_port, 
      RAM_2_90_port, RAM_2_89_port, RAM_2_88_port, RAM_2_87_port, RAM_2_86_port
      , RAM_2_85_port, RAM_2_84_port, RAM_2_83_port, RAM_2_82_port, 
      RAM_2_81_port, RAM_2_80_port, RAM_2_79_port, RAM_2_78_port, RAM_2_77_port
      , RAM_2_76_port, RAM_2_75_port, RAM_2_74_port, RAM_2_73_port, 
      RAM_2_72_port, RAM_2_71_port, RAM_2_70_port, RAM_2_69_port, RAM_2_68_port
      , RAM_2_67_port, RAM_2_66_port, RAM_2_65_port, RAM_2_64_port, 
      RAM_2_63_port, RAM_2_62_port, RAM_2_61_port, RAM_2_60_port, RAM_2_59_port
      , RAM_2_58_port, RAM_2_57_port, RAM_2_56_port, RAM_2_55_port, 
      RAM_2_54_port, RAM_2_53_port, RAM_2_52_port, RAM_2_51_port, RAM_2_50_port
      , RAM_2_49_port, RAM_2_48_port, RAM_2_47_port, RAM_2_46_port, 
      RAM_2_45_port, RAM_2_44_port, RAM_2_43_port, RAM_2_42_port, RAM_2_41_port
      , RAM_2_40_port, RAM_2_39_port, RAM_2_38_port, RAM_2_37_port, 
      RAM_2_36_port, RAM_2_35_port, RAM_2_34_port, RAM_2_33_port, RAM_2_32_port
      , RAM_2_31_port, RAM_2_30_port, RAM_2_29_port, RAM_2_28_port, 
      RAM_2_27_port, RAM_2_26_port, RAM_2_25_port, RAM_2_24_port, RAM_2_23_port
      , RAM_2_22_port, RAM_2_21_port, RAM_2_20_port, RAM_2_19_port, 
      RAM_2_18_port, RAM_2_17_port, RAM_2_16_port, RAM_2_15_port, RAM_2_14_port
      , RAM_2_13_port, RAM_2_12_port, RAM_2_11_port, RAM_2_10_port, 
      RAM_2_9_port, RAM_2_8_port, RAM_2_7_port, RAM_2_6_port, RAM_2_5_port, 
      RAM_2_4_port, RAM_2_3_port, RAM_2_2_port, RAM_2_1_port, RAM_2_0_port, 
      RAM_3_127_port, RAM_3_126_port, RAM_3_125_port, RAM_3_124_port, 
      RAM_3_123_port, RAM_3_122_port, RAM_3_121_port, RAM_3_120_port, 
      RAM_3_119_port, RAM_3_118_port, RAM_3_117_port, RAM_3_116_port, 
      RAM_3_115_port, RAM_3_114_port, RAM_3_113_port, RAM_3_112_port, 
      RAM_3_111_port, RAM_3_110_port, RAM_3_109_port, RAM_3_108_port, 
      RAM_3_107_port, RAM_3_106_port, RAM_3_105_port, RAM_3_104_port, 
      RAM_3_103_port, RAM_3_102_port, RAM_3_101_port, RAM_3_100_port, 
      RAM_3_99_port, RAM_3_98_port, RAM_3_97_port, RAM_3_96_port, RAM_3_95_port
      , RAM_3_94_port, RAM_3_93_port, RAM_3_92_port, RAM_3_91_port, 
      RAM_3_90_port, RAM_3_89_port, RAM_3_88_port, RAM_3_87_port, RAM_3_86_port
      , RAM_3_85_port, RAM_3_84_port, RAM_3_83_port, RAM_3_82_port, 
      RAM_3_81_port, RAM_3_80_port, RAM_3_79_port, RAM_3_78_port, RAM_3_77_port
      , RAM_3_76_port, RAM_3_75_port, RAM_3_74_port, RAM_3_73_port, 
      RAM_3_72_port, RAM_3_71_port, RAM_3_70_port, RAM_3_69_port, RAM_3_68_port
      , RAM_3_67_port, RAM_3_66_port, RAM_3_65_port, RAM_3_64_port, 
      RAM_3_63_port, RAM_3_62_port, RAM_3_61_port, RAM_3_60_port, RAM_3_59_port
      , RAM_3_58_port, RAM_3_57_port, RAM_3_56_port, RAM_3_55_port, 
      RAM_3_54_port, RAM_3_53_port, RAM_3_52_port, RAM_3_51_port, RAM_3_50_port
      , RAM_3_49_port, RAM_3_48_port, RAM_3_47_port, RAM_3_46_port, 
      RAM_3_45_port, RAM_3_44_port, RAM_3_43_port, RAM_3_42_port, RAM_3_41_port
      , RAM_3_40_port, RAM_3_39_port, RAM_3_38_port, RAM_3_37_port, 
      RAM_3_36_port, RAM_3_35_port, RAM_3_34_port, RAM_3_33_port, RAM_3_32_port
      , RAM_3_31_port, RAM_3_30_port, RAM_3_29_port, RAM_3_28_port, 
      RAM_3_27_port, RAM_3_26_port, RAM_3_25_port, RAM_3_24_port, RAM_3_23_port
      , RAM_3_22_port, RAM_3_21_port, RAM_3_20_port, RAM_3_19_port, 
      RAM_3_18_port, RAM_3_17_port, RAM_3_16_port, RAM_3_15_port, RAM_3_14_port
      , RAM_3_13_port, RAM_3_12_port, RAM_3_11_port, RAM_3_10_port, 
      RAM_3_9_port, RAM_3_8_port, RAM_3_7_port, RAM_3_6_port, RAM_3_5_port, 
      RAM_3_4_port, RAM_3_3_port, RAM_3_2_port, RAM_3_1_port, RAM_3_0_port, 
      RAM_4_127_port, RAM_4_126_port, RAM_4_125_port, RAM_4_124_port, 
      RAM_4_123_port, RAM_4_122_port, RAM_4_121_port, RAM_4_120_port, 
      RAM_4_119_port, RAM_4_118_port, RAM_4_117_port, RAM_4_116_port, 
      RAM_4_115_port, RAM_4_114_port, RAM_4_113_port, RAM_4_112_port, 
      RAM_4_111_port, RAM_4_110_port, RAM_4_109_port, RAM_4_108_port, 
      RAM_4_107_port, RAM_4_106_port, RAM_4_105_port, RAM_4_104_port, 
      RAM_4_103_port, RAM_4_102_port, RAM_4_101_port, RAM_4_100_port, 
      RAM_4_99_port, RAM_4_98_port, RAM_4_97_port, RAM_4_96_port, RAM_4_95_port
      , RAM_4_94_port, RAM_4_93_port, RAM_4_92_port, RAM_4_91_port, 
      RAM_4_90_port, RAM_4_89_port, RAM_4_88_port, RAM_4_87_port, RAM_4_86_port
      , RAM_4_85_port, RAM_4_84_port, RAM_4_83_port, RAM_4_82_port, 
      RAM_4_81_port, RAM_4_80_port, RAM_4_79_port, RAM_4_78_port, RAM_4_77_port
      , RAM_4_76_port, RAM_4_75_port, RAM_4_74_port, RAM_4_73_port, 
      RAM_4_72_port, RAM_4_71_port, RAM_4_70_port, RAM_4_69_port, RAM_4_68_port
      , RAM_4_67_port, RAM_4_66_port, RAM_4_65_port, RAM_4_64_port, 
      RAM_4_63_port, RAM_4_62_port, RAM_4_61_port, RAM_4_60_port, RAM_4_59_port
      , RAM_4_58_port, RAM_4_57_port, RAM_4_56_port, RAM_4_55_port, 
      RAM_4_54_port, RAM_4_53_port, RAM_4_52_port, RAM_4_51_port, RAM_4_50_port
      , RAM_4_49_port, RAM_4_48_port, RAM_4_47_port, RAM_4_46_port, 
      RAM_4_45_port, RAM_4_44_port, RAM_4_43_port, RAM_4_42_port, RAM_4_41_port
      , RAM_4_40_port, RAM_4_39_port, RAM_4_38_port, RAM_4_37_port, 
      RAM_4_36_port, RAM_4_35_port, RAM_4_34_port, RAM_4_33_port, RAM_4_32_port
      , RAM_4_31_port, RAM_4_30_port, RAM_4_29_port, RAM_4_28_port, 
      RAM_4_27_port, RAM_4_26_port, RAM_4_25_port, RAM_4_24_port, RAM_4_23_port
      , RAM_4_22_port, RAM_4_21_port, RAM_4_20_port, RAM_4_19_port, 
      RAM_4_18_port, RAM_4_17_port, RAM_4_16_port, RAM_4_15_port, RAM_4_14_port
      , RAM_4_13_port, RAM_4_12_port, RAM_4_11_port, RAM_4_10_port, 
      RAM_4_9_port, RAM_4_8_port, RAM_4_7_port, RAM_4_6_port, RAM_4_5_port, 
      RAM_4_4_port, RAM_4_3_port, RAM_4_2_port, RAM_4_1_port, RAM_4_0_port, 
      RAM_5_127_port, RAM_5_126_port, RAM_5_125_port, RAM_5_124_port, 
      RAM_5_123_port, RAM_5_122_port, RAM_5_121_port, RAM_5_120_port, 
      RAM_5_119_port, RAM_5_118_port, RAM_5_117_port, RAM_5_116_port, 
      RAM_5_115_port, RAM_5_114_port, RAM_5_113_port, RAM_5_112_port, 
      RAM_5_111_port, RAM_5_110_port, RAM_5_109_port, RAM_5_108_port, 
      RAM_5_107_port, RAM_5_106_port, RAM_5_105_port, RAM_5_104_port, 
      RAM_5_103_port, RAM_5_102_port, RAM_5_101_port, RAM_5_100_port, 
      RAM_5_99_port, RAM_5_98_port, RAM_5_97_port, RAM_5_96_port, RAM_5_95_port
      , RAM_5_94_port, RAM_5_93_port, RAM_5_92_port, RAM_5_91_port, 
      RAM_5_90_port, RAM_5_89_port, RAM_5_88_port, RAM_5_87_port, RAM_5_86_port
      , RAM_5_85_port, RAM_5_84_port, RAM_5_83_port, RAM_5_82_port, 
      RAM_5_81_port, RAM_5_80_port, RAM_5_79_port, RAM_5_78_port, RAM_5_77_port
      , RAM_5_76_port, RAM_5_75_port, RAM_5_74_port, RAM_5_73_port, 
      RAM_5_72_port, RAM_5_71_port, RAM_5_70_port, RAM_5_69_port, RAM_5_68_port
      , RAM_5_67_port, RAM_5_66_port, RAM_5_65_port, RAM_5_64_port, 
      RAM_5_63_port, RAM_5_62_port, RAM_5_61_port, RAM_5_60_port, RAM_5_59_port
      , RAM_5_58_port, RAM_5_57_port, RAM_5_56_port, RAM_5_55_port, 
      RAM_5_54_port, RAM_5_53_port, RAM_5_52_port, RAM_5_51_port, RAM_5_50_port
      , RAM_5_49_port, RAM_5_48_port, RAM_5_47_port, RAM_5_46_port, 
      RAM_5_45_port, RAM_5_44_port, RAM_5_43_port, RAM_5_42_port, RAM_5_41_port
      , RAM_5_40_port, RAM_5_39_port, RAM_5_38_port, RAM_5_37_port, 
      RAM_5_36_port, RAM_5_35_port, RAM_5_34_port, RAM_5_33_port, RAM_5_32_port
      , RAM_5_31_port, RAM_5_30_port, RAM_5_29_port, RAM_5_28_port, 
      RAM_5_27_port, RAM_5_26_port, RAM_5_25_port, RAM_5_24_port, RAM_5_23_port
      , RAM_5_22_port, RAM_5_21_port, RAM_5_20_port, RAM_5_19_port, 
      RAM_5_18_port, RAM_5_17_port, RAM_5_16_port, RAM_5_15_port, RAM_5_14_port
      , RAM_5_13_port, RAM_5_12_port, RAM_5_11_port, RAM_5_10_port, 
      RAM_5_9_port, RAM_5_8_port, RAM_5_7_port, RAM_5_6_port, RAM_5_5_port, 
      RAM_5_4_port, RAM_5_3_port, RAM_5_2_port, RAM_5_1_port, RAM_5_0_port, 
      RAM_6_127_port, RAM_6_126_port, RAM_6_125_port, RAM_6_124_port, 
      RAM_6_123_port, RAM_6_122_port, RAM_6_121_port, RAM_6_120_port, 
      RAM_6_119_port, RAM_6_118_port, RAM_6_117_port, RAM_6_116_port, 
      RAM_6_115_port, RAM_6_114_port, RAM_6_113_port, RAM_6_112_port, 
      RAM_6_111_port, RAM_6_110_port, RAM_6_109_port, RAM_6_108_port, 
      RAM_6_107_port, RAM_6_106_port, RAM_6_105_port, RAM_6_104_port, 
      RAM_6_103_port, RAM_6_102_port, RAM_6_101_port, RAM_6_100_port, 
      RAM_6_99_port, RAM_6_98_port, RAM_6_97_port, RAM_6_96_port, RAM_6_95_port
      , RAM_6_94_port, RAM_6_93_port, RAM_6_92_port, RAM_6_91_port, 
      RAM_6_90_port, RAM_6_89_port, RAM_6_88_port, RAM_6_87_port, RAM_6_86_port
      , RAM_6_85_port, RAM_6_84_port, RAM_6_83_port, RAM_6_82_port, 
      RAM_6_81_port, RAM_6_80_port, RAM_6_79_port, RAM_6_78_port, RAM_6_77_port
      , RAM_6_76_port, RAM_6_75_port, RAM_6_74_port, RAM_6_73_port, 
      RAM_6_72_port, RAM_6_71_port, RAM_6_70_port, RAM_6_69_port, RAM_6_68_port
      , RAM_6_67_port, RAM_6_66_port, RAM_6_65_port, RAM_6_64_port, 
      RAM_6_63_port, RAM_6_62_port, RAM_6_61_port, RAM_6_60_port, RAM_6_59_port
      , RAM_6_58_port, RAM_6_57_port, RAM_6_56_port, RAM_6_55_port, 
      RAM_6_54_port, RAM_6_53_port, RAM_6_52_port, RAM_6_51_port, RAM_6_50_port
      , RAM_6_49_port, RAM_6_48_port, RAM_6_47_port, RAM_6_46_port, 
      RAM_6_45_port, RAM_6_44_port, RAM_6_43_port, RAM_6_42_port, RAM_6_41_port
      , RAM_6_40_port, RAM_6_39_port, RAM_6_38_port, RAM_6_37_port, 
      RAM_6_36_port, RAM_6_35_port, RAM_6_34_port, RAM_6_33_port, RAM_6_32_port
      , RAM_6_31_port, RAM_6_30_port, RAM_6_29_port, RAM_6_28_port, 
      RAM_6_27_port, RAM_6_26_port, RAM_6_25_port, RAM_6_24_port, RAM_6_23_port
      , RAM_6_22_port, RAM_6_21_port, RAM_6_20_port, RAM_6_19_port, 
      RAM_6_18_port, RAM_6_17_port, RAM_6_16_port, RAM_6_15_port, RAM_6_14_port
      , RAM_6_13_port, RAM_6_12_port, RAM_6_11_port, RAM_6_10_port, 
      RAM_6_9_port, RAM_6_8_port, RAM_6_7_port, RAM_6_6_port, RAM_6_5_port, 
      RAM_6_4_port, RAM_6_3_port, RAM_6_2_port, RAM_6_1_port, RAM_6_0_port, 
      RAM_7_127_port, RAM_7_126_port, RAM_7_125_port, RAM_7_124_port, 
      RAM_7_123_port, RAM_7_122_port, RAM_7_121_port, RAM_7_120_port, 
      RAM_7_119_port, RAM_7_118_port, RAM_7_117_port, RAM_7_116_port, 
      RAM_7_115_port, RAM_7_114_port, RAM_7_113_port, RAM_7_112_port, 
      RAM_7_111_port, RAM_7_110_port, RAM_7_109_port, RAM_7_108_port, 
      RAM_7_107_port, RAM_7_106_port, RAM_7_105_port, RAM_7_104_port, 
      RAM_7_103_port, RAM_7_102_port, RAM_7_101_port, RAM_7_100_port, 
      RAM_7_99_port, RAM_7_98_port, RAM_7_97_port, RAM_7_96_port, RAM_7_95_port
      , RAM_7_94_port, RAM_7_93_port, RAM_7_92_port, RAM_7_91_port, 
      RAM_7_90_port, RAM_7_89_port, RAM_7_88_port, RAM_7_87_port, RAM_7_86_port
      , RAM_7_85_port, RAM_7_84_port, RAM_7_83_port, RAM_7_82_port, 
      RAM_7_81_port, RAM_7_80_port, RAM_7_79_port, RAM_7_78_port, RAM_7_77_port
      , RAM_7_76_port, RAM_7_75_port, RAM_7_74_port, RAM_7_73_port, 
      RAM_7_72_port, RAM_7_71_port, RAM_7_70_port, RAM_7_69_port, RAM_7_68_port
      , RAM_7_67_port, RAM_7_66_port, RAM_7_65_port, RAM_7_64_port, 
      RAM_7_63_port, RAM_7_62_port, RAM_7_61_port, RAM_7_60_port, RAM_7_59_port
      , RAM_7_58_port, RAM_7_57_port, RAM_7_56_port, RAM_7_55_port, 
      RAM_7_54_port, RAM_7_53_port, RAM_7_52_port, RAM_7_51_port, RAM_7_50_port
      , RAM_7_49_port, RAM_7_48_port, RAM_7_47_port, RAM_7_46_port, 
      RAM_7_45_port, RAM_7_44_port, RAM_7_43_port, RAM_7_42_port, RAM_7_41_port
      , RAM_7_40_port, RAM_7_39_port, RAM_7_38_port, RAM_7_37_port, 
      RAM_7_36_port, RAM_7_35_port, RAM_7_34_port, RAM_7_33_port, RAM_7_32_port
      , RAM_7_31_port, RAM_7_30_port, RAM_7_29_port, RAM_7_28_port, 
      RAM_7_27_port, RAM_7_26_port, RAM_7_25_port, RAM_7_24_port, RAM_7_23_port
      , RAM_7_22_port, RAM_7_21_port, RAM_7_20_port, RAM_7_19_port, 
      RAM_7_18_port, RAM_7_17_port, RAM_7_16_port, RAM_7_15_port, RAM_7_14_port
      , RAM_7_13_port, RAM_7_12_port, RAM_7_11_port, RAM_7_10_port, 
      RAM_7_9_port, RAM_7_8_port, RAM_7_7_port, RAM_7_6_port, RAM_7_5_port, 
      RAM_7_4_port, RAM_7_3_port, RAM_7_2_port, RAM_7_1_port, RAM_7_0_port, 
      RAM_8_127_port, RAM_8_126_port, RAM_8_125_port, RAM_8_124_port, 
      RAM_8_123_port, RAM_8_122_port, RAM_8_121_port, RAM_8_120_port, 
      RAM_8_119_port, RAM_8_118_port, RAM_8_117_port, RAM_8_116_port, 
      RAM_8_115_port, RAM_8_114_port, RAM_8_113_port, RAM_8_112_port, 
      RAM_8_111_port, RAM_8_110_port, RAM_8_109_port, RAM_8_108_port, 
      RAM_8_107_port, RAM_8_106_port, RAM_8_105_port, RAM_8_104_port, 
      RAM_8_103_port, RAM_8_102_port, RAM_8_101_port, RAM_8_100_port, 
      RAM_8_99_port, RAM_8_98_port, RAM_8_97_port, RAM_8_96_port, RAM_8_95_port
      , RAM_8_94_port, RAM_8_93_port, RAM_8_92_port, RAM_8_91_port, 
      RAM_8_90_port, RAM_8_89_port, RAM_8_88_port, RAM_8_87_port, RAM_8_86_port
      , RAM_8_85_port, RAM_8_84_port, RAM_8_83_port, RAM_8_82_port, 
      RAM_8_81_port, RAM_8_80_port, RAM_8_79_port, RAM_8_78_port, RAM_8_77_port
      , RAM_8_76_port, RAM_8_75_port, RAM_8_74_port, RAM_8_73_port, 
      RAM_8_72_port, RAM_8_71_port, RAM_8_70_port, RAM_8_69_port, RAM_8_68_port
      , RAM_8_67_port, RAM_8_66_port, RAM_8_65_port, RAM_8_64_port, 
      RAM_8_63_port, RAM_8_62_port, RAM_8_61_port, RAM_8_60_port, RAM_8_59_port
      , RAM_8_58_port, RAM_8_57_port, RAM_8_56_port, RAM_8_55_port, 
      RAM_8_54_port, RAM_8_53_port, RAM_8_52_port, RAM_8_51_port, RAM_8_50_port
      , RAM_8_49_port, RAM_8_48_port, RAM_8_47_port, RAM_8_46_port, 
      RAM_8_45_port, RAM_8_44_port, RAM_8_43_port, RAM_8_42_port, RAM_8_41_port
      , RAM_8_40_port, RAM_8_39_port, RAM_8_38_port, RAM_8_37_port, 
      RAM_8_36_port, RAM_8_35_port, RAM_8_34_port, RAM_8_33_port, RAM_8_32_port
      , RAM_8_31_port, RAM_8_30_port, RAM_8_29_port, RAM_8_28_port, 
      RAM_8_27_port, RAM_8_26_port, RAM_8_25_port, RAM_8_24_port, RAM_8_23_port
      , RAM_8_22_port, RAM_8_21_port, RAM_8_20_port, RAM_8_19_port, 
      RAM_8_18_port, RAM_8_17_port, RAM_8_16_port, RAM_8_15_port, RAM_8_14_port
      , RAM_8_13_port, RAM_8_12_port, RAM_8_11_port, RAM_8_10_port, 
      RAM_8_9_port, RAM_8_8_port, RAM_8_7_port, RAM_8_6_port, RAM_8_5_port, 
      RAM_8_4_port, RAM_8_3_port, RAM_8_2_port, RAM_8_1_port, RAM_8_0_port, 
      RAM_9_127_port, RAM_9_126_port, RAM_9_125_port, RAM_9_124_port, 
      RAM_9_123_port, RAM_9_122_port, RAM_9_121_port, RAM_9_120_port, 
      RAM_9_119_port, RAM_9_118_port, RAM_9_117_port, RAM_9_116_port, 
      RAM_9_115_port, RAM_9_114_port, RAM_9_113_port, RAM_9_112_port, 
      RAM_9_111_port, RAM_9_110_port, RAM_9_109_port, RAM_9_108_port, 
      RAM_9_107_port, RAM_9_106_port, RAM_9_105_port, RAM_9_104_port, 
      RAM_9_103_port, RAM_9_102_port, RAM_9_101_port, RAM_9_100_port, 
      RAM_9_99_port, RAM_9_98_port, RAM_9_97_port, RAM_9_96_port, RAM_9_95_port
      , RAM_9_94_port, RAM_9_93_port, RAM_9_92_port, RAM_9_91_port, 
      RAM_9_90_port, RAM_9_89_port, RAM_9_88_port, RAM_9_87_port, RAM_9_86_port
      , RAM_9_85_port, RAM_9_84_port, RAM_9_83_port, RAM_9_82_port, 
      RAM_9_81_port, RAM_9_80_port, RAM_9_79_port, RAM_9_78_port, RAM_9_77_port
      , RAM_9_76_port, RAM_9_75_port, RAM_9_74_port, RAM_9_73_port, 
      RAM_9_72_port, RAM_9_71_port, RAM_9_70_port, RAM_9_69_port, RAM_9_68_port
      , RAM_9_67_port, RAM_9_66_port, RAM_9_65_port, RAM_9_64_port, 
      RAM_9_63_port, RAM_9_62_port, RAM_9_61_port, RAM_9_60_port, RAM_9_59_port
      , RAM_9_58_port, RAM_9_57_port, RAM_9_56_port, RAM_9_55_port, 
      RAM_9_54_port, RAM_9_53_port, RAM_9_52_port, RAM_9_51_port, RAM_9_50_port
      , RAM_9_49_port, RAM_9_48_port, RAM_9_47_port, RAM_9_46_port, 
      RAM_9_45_port, RAM_9_44_port, RAM_9_43_port, RAM_9_42_port, RAM_9_41_port
      , RAM_9_40_port, RAM_9_39_port, RAM_9_38_port, RAM_9_37_port, 
      RAM_9_36_port, RAM_9_35_port, RAM_9_34_port, RAM_9_33_port, RAM_9_32_port
      , RAM_9_31_port, RAM_9_30_port, RAM_9_29_port, RAM_9_28_port, 
      RAM_9_27_port, RAM_9_26_port, RAM_9_25_port, RAM_9_24_port, RAM_9_23_port
      , RAM_9_22_port, RAM_9_21_port, RAM_9_20_port, RAM_9_19_port, 
      RAM_9_18_port, RAM_9_17_port, RAM_9_16_port, RAM_9_15_port, RAM_9_14_port
      , RAM_9_13_port, RAM_9_12_port, RAM_9_11_port, RAM_9_10_port, 
      RAM_9_9_port, RAM_9_8_port, RAM_9_7_port, RAM_9_6_port, RAM_9_5_port, 
      RAM_9_4_port, RAM_9_3_port, RAM_9_2_port, RAM_9_1_port, RAM_9_0_port, 
      RAM_10_127_port, RAM_10_126_port, RAM_10_125_port, RAM_10_124_port, 
      RAM_10_123_port, RAM_10_122_port, RAM_10_121_port, RAM_10_120_port, 
      RAM_10_119_port, RAM_10_118_port, RAM_10_117_port, RAM_10_116_port, 
      RAM_10_115_port, RAM_10_114_port, RAM_10_113_port, RAM_10_112_port, 
      RAM_10_111_port, RAM_10_110_port, RAM_10_109_port, RAM_10_108_port, 
      RAM_10_107_port, RAM_10_106_port, RAM_10_105_port, RAM_10_104_port, 
      RAM_10_103_port, RAM_10_102_port, RAM_10_101_port, RAM_10_100_port, 
      RAM_10_99_port, RAM_10_98_port, RAM_10_97_port, RAM_10_96_port, 
      RAM_10_95_port, RAM_10_94_port, RAM_10_93_port, RAM_10_92_port, 
      RAM_10_91_port, RAM_10_90_port, RAM_10_89_port, RAM_10_88_port, 
      RAM_10_87_port, RAM_10_86_port, RAM_10_85_port, RAM_10_84_port, 
      RAM_10_83_port, RAM_10_82_port, RAM_10_81_port, RAM_10_80_port, 
      RAM_10_79_port, RAM_10_78_port, RAM_10_77_port, RAM_10_76_port, 
      RAM_10_75_port, RAM_10_74_port, RAM_10_73_port, RAM_10_72_port, 
      RAM_10_71_port, RAM_10_70_port, RAM_10_69_port, RAM_10_68_port, 
      RAM_10_67_port, RAM_10_66_port, RAM_10_65_port, RAM_10_64_port, 
      RAM_10_63_port, RAM_10_62_port, RAM_10_61_port, RAM_10_60_port, 
      RAM_10_59_port, RAM_10_58_port, RAM_10_57_port, RAM_10_56_port, 
      RAM_10_55_port, RAM_10_54_port, RAM_10_53_port, RAM_10_52_port, 
      RAM_10_51_port, RAM_10_50_port, RAM_10_49_port, RAM_10_48_port, 
      RAM_10_47_port, RAM_10_46_port, RAM_10_45_port, RAM_10_44_port, 
      RAM_10_43_port, RAM_10_42_port, RAM_10_41_port, RAM_10_40_port, 
      RAM_10_39_port, RAM_10_38_port, RAM_10_37_port, RAM_10_36_port, 
      RAM_10_35_port, RAM_10_34_port, RAM_10_33_port, RAM_10_32_port, 
      RAM_10_31_port, RAM_10_30_port, RAM_10_29_port, RAM_10_28_port, 
      RAM_10_27_port, RAM_10_26_port, RAM_10_25_port, RAM_10_24_port, 
      RAM_10_23_port, RAM_10_22_port, RAM_10_21_port, RAM_10_20_port, 
      RAM_10_19_port, RAM_10_18_port, RAM_10_17_port, RAM_10_16_port, 
      RAM_10_15_port, RAM_10_14_port, RAM_10_13_port, RAM_10_12_port, 
      RAM_10_11_port, RAM_10_10_port, RAM_10_9_port, RAM_10_8_port, 
      RAM_10_7_port, RAM_10_6_port, RAM_10_5_port, RAM_10_4_port, RAM_10_3_port
      , RAM_10_2_port, RAM_10_1_port, RAM_10_0_port, RAM_11_127_port, 
      RAM_11_126_port, RAM_11_125_port, RAM_11_124_port, RAM_11_123_port, 
      RAM_11_122_port, RAM_11_121_port, RAM_11_120_port, RAM_11_119_port, 
      RAM_11_118_port, RAM_11_117_port, RAM_11_116_port, RAM_11_115_port, 
      RAM_11_114_port, RAM_11_113_port, RAM_11_112_port, RAM_11_111_port, 
      RAM_11_110_port, RAM_11_109_port, RAM_11_108_port, RAM_11_107_port, 
      RAM_11_106_port, RAM_11_105_port, RAM_11_104_port, RAM_11_103_port, 
      RAM_11_102_port, RAM_11_101_port, RAM_11_100_port, RAM_11_99_port, 
      RAM_11_98_port, RAM_11_97_port, RAM_11_96_port, RAM_11_95_port, 
      RAM_11_94_port, RAM_11_93_port, RAM_11_92_port, RAM_11_91_port, 
      RAM_11_90_port, RAM_11_89_port, RAM_11_88_port, RAM_11_87_port, 
      RAM_11_86_port, RAM_11_85_port, RAM_11_84_port, RAM_11_83_port, 
      RAM_11_82_port, RAM_11_81_port, RAM_11_80_port, RAM_11_79_port, 
      RAM_11_78_port, RAM_11_77_port, RAM_11_76_port, RAM_11_75_port, 
      RAM_11_74_port, RAM_11_73_port, RAM_11_72_port, RAM_11_71_port, 
      RAM_11_70_port, RAM_11_69_port, RAM_11_68_port, RAM_11_67_port, 
      RAM_11_66_port, RAM_11_65_port, RAM_11_64_port, RAM_11_63_port, 
      RAM_11_62_port, RAM_11_61_port, RAM_11_60_port, RAM_11_59_port, 
      RAM_11_58_port, RAM_11_57_port, RAM_11_56_port, RAM_11_55_port, 
      RAM_11_54_port, RAM_11_53_port, RAM_11_52_port, RAM_11_51_port, 
      RAM_11_50_port, RAM_11_49_port, RAM_11_48_port, RAM_11_47_port, 
      RAM_11_46_port, RAM_11_45_port, RAM_11_44_port, RAM_11_43_port, 
      RAM_11_42_port, RAM_11_41_port, RAM_11_40_port, RAM_11_39_port, 
      RAM_11_38_port, RAM_11_37_port, RAM_11_36_port, RAM_11_35_port, 
      RAM_11_34_port, RAM_11_33_port, RAM_11_32_port, RAM_11_31_port, 
      RAM_11_30_port, RAM_11_29_port, RAM_11_28_port, RAM_11_27_port, 
      RAM_11_26_port, RAM_11_25_port, RAM_11_24_port, RAM_11_23_port, 
      RAM_11_22_port, RAM_11_21_port, RAM_11_20_port, RAM_11_19_port, 
      RAM_11_18_port, RAM_11_17_port, RAM_11_16_port, RAM_11_15_port, 
      RAM_11_14_port, RAM_11_13_port, RAM_11_12_port, RAM_11_11_port, 
      RAM_11_10_port, RAM_11_9_port, RAM_11_8_port, RAM_11_7_port, 
      RAM_11_6_port, RAM_11_5_port, RAM_11_4_port, RAM_11_3_port, RAM_11_2_port
      , RAM_11_1_port, RAM_11_0_port, RAM_12_127_port, RAM_12_126_port, 
      RAM_12_125_port, RAM_12_124_port, RAM_12_123_port, RAM_12_122_port, 
      RAM_12_121_port, RAM_12_120_port, RAM_12_119_port, RAM_12_118_port, 
      RAM_12_117_port, RAM_12_116_port, RAM_12_115_port, RAM_12_114_port, 
      RAM_12_113_port, RAM_12_112_port, RAM_12_111_port, RAM_12_110_port, 
      RAM_12_109_port, RAM_12_108_port, RAM_12_107_port, RAM_12_106_port, 
      RAM_12_105_port, RAM_12_104_port, RAM_12_103_port, RAM_12_102_port, 
      RAM_12_101_port, RAM_12_100_port, RAM_12_99_port, RAM_12_98_port, 
      RAM_12_97_port, RAM_12_96_port, RAM_12_95_port, RAM_12_94_port, 
      RAM_12_93_port, RAM_12_92_port, RAM_12_91_port, RAM_12_90_port, 
      RAM_12_89_port, RAM_12_88_port, RAM_12_87_port, RAM_12_86_port, 
      RAM_12_85_port, RAM_12_84_port, RAM_12_83_port, RAM_12_82_port, 
      RAM_12_81_port, RAM_12_80_port, RAM_12_79_port, RAM_12_78_port, 
      RAM_12_77_port, RAM_12_76_port, RAM_12_75_port, RAM_12_74_port, 
      RAM_12_73_port, RAM_12_72_port, RAM_12_71_port, RAM_12_70_port, 
      RAM_12_69_port, RAM_12_68_port, RAM_12_67_port, RAM_12_66_port, 
      RAM_12_65_port, RAM_12_64_port, RAM_12_63_port, RAM_12_62_port, 
      RAM_12_61_port, RAM_12_60_port, RAM_12_59_port, RAM_12_58_port, 
      RAM_12_57_port, RAM_12_56_port, RAM_12_55_port, RAM_12_54_port, 
      RAM_12_53_port, RAM_12_52_port, RAM_12_51_port, RAM_12_50_port, 
      RAM_12_49_port, RAM_12_48_port, RAM_12_47_port, RAM_12_46_port, 
      RAM_12_45_port, RAM_12_44_port, RAM_12_43_port, RAM_12_42_port, 
      RAM_12_41_port, RAM_12_40_port, RAM_12_39_port, RAM_12_38_port, 
      RAM_12_37_port, RAM_12_36_port, RAM_12_35_port, RAM_12_34_port, 
      RAM_12_33_port, RAM_12_32_port, RAM_12_31_port, RAM_12_30_port, 
      RAM_12_29_port, RAM_12_28_port, RAM_12_27_port, RAM_12_26_port, 
      RAM_12_25_port, RAM_12_24_port, RAM_12_23_port, RAM_12_22_port, 
      RAM_12_21_port, RAM_12_20_port, RAM_12_19_port, RAM_12_18_port, 
      RAM_12_17_port, RAM_12_16_port, RAM_12_15_port, RAM_12_14_port, 
      RAM_12_13_port, RAM_12_12_port, RAM_12_11_port, RAM_12_10_port, 
      RAM_12_9_port, RAM_12_8_port, RAM_12_7_port, RAM_12_6_port, RAM_12_5_port
      , RAM_12_4_port, RAM_12_3_port, RAM_12_2_port, RAM_12_1_port, 
      RAM_12_0_port, RAM_13_127_port, RAM_13_126_port, RAM_13_125_port, 
      RAM_13_124_port, RAM_13_123_port, RAM_13_122_port, RAM_13_121_port, 
      RAM_13_120_port, RAM_13_119_port, RAM_13_118_port, RAM_13_117_port, 
      RAM_13_116_port, RAM_13_115_port, RAM_13_114_port, RAM_13_113_port, 
      RAM_13_112_port, RAM_13_111_port, RAM_13_110_port, RAM_13_109_port, 
      RAM_13_108_port, RAM_13_107_port, RAM_13_106_port, RAM_13_105_port, 
      RAM_13_104_port, RAM_13_103_port, RAM_13_102_port, RAM_13_101_port, 
      RAM_13_100_port, RAM_13_99_port, RAM_13_98_port, RAM_13_97_port, 
      RAM_13_96_port, RAM_13_95_port, RAM_13_94_port, RAM_13_93_port, 
      RAM_13_92_port, RAM_13_91_port, RAM_13_90_port, RAM_13_89_port, 
      RAM_13_88_port, RAM_13_87_port, RAM_13_86_port, RAM_13_85_port, 
      RAM_13_84_port, RAM_13_83_port, RAM_13_82_port, RAM_13_81_port, 
      RAM_13_80_port, RAM_13_79_port, RAM_13_78_port, RAM_13_77_port, 
      RAM_13_76_port, RAM_13_75_port, RAM_13_74_port, RAM_13_73_port, 
      RAM_13_72_port, RAM_13_71_port, RAM_13_70_port, RAM_13_69_port, 
      RAM_13_68_port, RAM_13_67_port, RAM_13_66_port, RAM_13_65_port, 
      RAM_13_64_port, RAM_13_63_port, RAM_13_62_port, RAM_13_61_port, 
      RAM_13_60_port, RAM_13_59_port, RAM_13_58_port, RAM_13_57_port, 
      RAM_13_56_port, RAM_13_55_port, RAM_13_54_port, RAM_13_53_port, 
      RAM_13_52_port, RAM_13_51_port, RAM_13_50_port, RAM_13_49_port, 
      RAM_13_48_port, RAM_13_47_port, RAM_13_46_port, RAM_13_45_port, 
      RAM_13_44_port, RAM_13_43_port, RAM_13_42_port, RAM_13_41_port, 
      RAM_13_40_port, RAM_13_39_port, RAM_13_38_port, RAM_13_37_port, 
      RAM_13_36_port, RAM_13_35_port, RAM_13_34_port, RAM_13_33_port, 
      RAM_13_32_port, RAM_13_31_port, RAM_13_30_port, RAM_13_29_port, 
      RAM_13_28_port, RAM_13_27_port, RAM_13_26_port, RAM_13_25_port, 
      RAM_13_24_port, RAM_13_23_port, RAM_13_22_port, RAM_13_21_port, 
      RAM_13_20_port, RAM_13_19_port, RAM_13_18_port, RAM_13_17_port, 
      RAM_13_16_port, RAM_13_15_port, RAM_13_14_port, RAM_13_13_port, 
      RAM_13_12_port, RAM_13_11_port, RAM_13_10_port, RAM_13_9_port, 
      RAM_13_8_port, RAM_13_7_port, RAM_13_6_port, RAM_13_5_port, RAM_13_4_port
      , RAM_13_3_port, RAM_13_2_port, RAM_13_1_port, RAM_13_0_port, 
      RAM_14_127_port, RAM_14_126_port, RAM_14_125_port, RAM_14_124_port, 
      RAM_14_123_port, RAM_14_122_port, RAM_14_121_port, RAM_14_120_port, 
      RAM_14_119_port, RAM_14_118_port, RAM_14_117_port, RAM_14_116_port, 
      RAM_14_115_port, RAM_14_114_port, RAM_14_113_port, RAM_14_112_port, 
      RAM_14_111_port, RAM_14_110_port, RAM_14_109_port, RAM_14_108_port, 
      RAM_14_107_port, RAM_14_106_port, RAM_14_105_port, RAM_14_104_port, 
      RAM_14_103_port, RAM_14_102_port, RAM_14_101_port, RAM_14_100_port, 
      RAM_14_99_port, RAM_14_98_port, RAM_14_97_port, RAM_14_96_port, 
      RAM_14_95_port, RAM_14_94_port, RAM_14_93_port, RAM_14_92_port, 
      RAM_14_91_port, RAM_14_90_port, RAM_14_89_port, RAM_14_88_port, 
      RAM_14_87_port, RAM_14_86_port, RAM_14_85_port, RAM_14_84_port, 
      RAM_14_83_port, RAM_14_82_port, RAM_14_81_port, RAM_14_80_port, 
      RAM_14_79_port, RAM_14_78_port, RAM_14_77_port, RAM_14_76_port, 
      RAM_14_75_port, RAM_14_74_port, RAM_14_73_port, RAM_14_72_port, 
      RAM_14_71_port, RAM_14_70_port, RAM_14_69_port, RAM_14_68_port, 
      RAM_14_67_port, RAM_14_66_port, RAM_14_65_port, RAM_14_64_port, 
      RAM_14_63_port, RAM_14_62_port, RAM_14_61_port, RAM_14_60_port, 
      RAM_14_59_port, RAM_14_58_port, RAM_14_57_port, RAM_14_56_port, 
      RAM_14_55_port, RAM_14_54_port, RAM_14_53_port, RAM_14_52_port, 
      RAM_14_51_port, RAM_14_50_port, RAM_14_49_port, RAM_14_48_port, 
      RAM_14_47_port, RAM_14_46_port, RAM_14_45_port, RAM_14_44_port, 
      RAM_14_43_port, RAM_14_42_port, RAM_14_41_port, RAM_14_40_port, 
      RAM_14_39_port, RAM_14_38_port, RAM_14_37_port, RAM_14_36_port, 
      RAM_14_35_port, RAM_14_34_port, RAM_14_33_port, RAM_14_32_port, 
      RAM_14_31_port, RAM_14_30_port, RAM_14_29_port, RAM_14_28_port, 
      RAM_14_27_port, RAM_14_26_port, RAM_14_25_port, RAM_14_24_port, 
      RAM_14_23_port, RAM_14_22_port, RAM_14_21_port, RAM_14_20_port, 
      RAM_14_19_port, RAM_14_18_port, RAM_14_17_port, RAM_14_16_port, 
      RAM_14_15_port, RAM_14_14_port, RAM_14_13_port, RAM_14_12_port, 
      RAM_14_11_port, RAM_14_10_port, RAM_14_9_port, RAM_14_8_port, 
      RAM_14_7_port, RAM_14_6_port, RAM_14_5_port, RAM_14_4_port, RAM_14_3_port
      , RAM_14_2_port, RAM_14_1_port, RAM_14_0_port, RAM_15_127_port, 
      RAM_15_126_port, RAM_15_125_port, RAM_15_124_port, RAM_15_123_port, 
      RAM_15_122_port, RAM_15_121_port, RAM_15_120_port, RAM_15_119_port, 
      RAM_15_118_port, RAM_15_117_port, RAM_15_116_port, RAM_15_115_port, 
      RAM_15_114_port, RAM_15_113_port, RAM_15_112_port, RAM_15_111_port, 
      RAM_15_110_port, RAM_15_109_port, RAM_15_108_port, RAM_15_107_port, 
      RAM_15_106_port, RAM_15_105_port, RAM_15_104_port, RAM_15_103_port, 
      RAM_15_102_port, RAM_15_101_port, RAM_15_100_port, RAM_15_99_port, 
      RAM_15_98_port, RAM_15_97_port, RAM_15_96_port, RAM_15_95_port, 
      RAM_15_94_port, RAM_15_93_port, RAM_15_92_port, RAM_15_91_port, 
      RAM_15_90_port, RAM_15_89_port, RAM_15_88_port, RAM_15_87_port, 
      RAM_15_86_port, RAM_15_85_port, RAM_15_84_port, RAM_15_83_port, 
      RAM_15_82_port, RAM_15_81_port, RAM_15_80_port, RAM_15_79_port, 
      RAM_15_78_port, RAM_15_77_port, RAM_15_76_port, RAM_15_75_port, 
      RAM_15_74_port, RAM_15_73_port, RAM_15_72_port, RAM_15_71_port, 
      RAM_15_70_port, RAM_15_69_port, RAM_15_68_port, RAM_15_67_port, 
      RAM_15_66_port, RAM_15_65_port, RAM_15_64_port, RAM_15_63_port, 
      RAM_15_62_port, RAM_15_61_port, RAM_15_60_port, RAM_15_59_port, 
      RAM_15_58_port, RAM_15_57_port, RAM_15_56_port, RAM_15_55_port, 
      RAM_15_54_port, RAM_15_53_port, RAM_15_52_port, RAM_15_51_port, 
      RAM_15_50_port, RAM_15_49_port, RAM_15_48_port, RAM_15_47_port, 
      RAM_15_46_port, RAM_15_45_port, RAM_15_44_port, RAM_15_43_port, 
      RAM_15_42_port, RAM_15_41_port, RAM_15_40_port, RAM_15_39_port, 
      RAM_15_38_port, RAM_15_37_port, RAM_15_36_port, RAM_15_35_port, 
      RAM_15_34_port, RAM_15_33_port, RAM_15_32_port, RAM_15_31_port, 
      RAM_15_30_port, RAM_15_29_port, RAM_15_28_port, RAM_15_27_port, 
      RAM_15_26_port, RAM_15_25_port, RAM_15_24_port, RAM_15_23_port, 
      RAM_15_22_port, RAM_15_21_port, RAM_15_20_port, RAM_15_19_port, 
      RAM_15_18_port, RAM_15_17_port, RAM_15_16_port, RAM_15_15_port, 
      RAM_15_14_port, RAM_15_13_port, RAM_15_12_port, RAM_15_11_port, 
      RAM_15_10_port, RAM_15_9_port, RAM_15_8_port, RAM_15_7_port, 
      RAM_15_6_port, RAM_15_5_port, RAM_15_4_port, RAM_15_3_port, RAM_15_2_port
      , RAM_15_1_port, RAM_15_0_port, n21, n22, n23, n24, n25, n26, n27, n28, 
      n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43
      , n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, 
      n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72
      , n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, 
      n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, 
      n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, 
      n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, 
      n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, 
      n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, 
      n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, 
      n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, 
      n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, 
      n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, 
      n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, 
      n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, 
      n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, 
      n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, 
      n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, 
      n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, 
      n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, 
      n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, 
      n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, 
      n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, 
      n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, 
      n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, 
      n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, 
      n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, 
      n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, 
      n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, 
      n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, 
      n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, 
      n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, 
      n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, 
      n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, 
      n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, 
      n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, 
      n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, 
      n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, 
      n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, 
      n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, 
      n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, 
      n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, 
      n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, 
      n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, 
      n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, 
      n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, 
      n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, 
      n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, 
      n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, 
      n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, 
      n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, 
      n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, 
      n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, 
      n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, 
      n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, 
      n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, 
      n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, 
      n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, 
      n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, 
      n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, 
      n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, 
      n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, 
      n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, 
      n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, 
      n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, 
      n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, 
      n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, 
      n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, 
      n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, 
      n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, 
      n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, 
      n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, 
      n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, 
      n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, 
      n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, 
      n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, 
      n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, 
      n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, 
      n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, 
      n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, 
      n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, 
      n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, 
      n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, 
      n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, 
      n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, 
      n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, 
      n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, 
      n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, 
      n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, 
      n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, 
      n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, 
      n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, 
      n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, 
      n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, 
      n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, 
      n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, 
      n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, 
      n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, 
      n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, 
      n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, 
      n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, 
      n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, 
      n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, 
      n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, 
      n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, 
      n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, 
      n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, 
      n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, 
      n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, 
      n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, 
      n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, 
      n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, 
      n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, 
      n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, 
      n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, 
      n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, 
      n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, 
      n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, 
      n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, 
      n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, 
      n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, 
      n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, 
      n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, 
      n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, 
      n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, 
      n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, 
      n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, 
      n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, 
      n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, 
      n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, 
      n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, 
      n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, 
      n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, 
      n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, 
      n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, 
      n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, 
      n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, 
      n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, 
      n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, 
      n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, 
      n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, 
      n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, 
      n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, 
      n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, 
      n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, 
      n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, 
      n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, 
      n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, 
      n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, 
      n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, 
      n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, 
      n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, 
      n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, 
      n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, 
      n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, 
      n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, 
      n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, 
      n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, 
      n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, 
      n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, 
      n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, 
      n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, 
      n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, 
      n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, 
      n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, 
      n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, 
      n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, 
      n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, 
      n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, 
      n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, 
      n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, 
      n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, 
      n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, 
      n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, 
      n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, 
      n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, 
      n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, 
      n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, 
      n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, 
      n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, 
      n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, 
      n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, 
      n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, 
      n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, 
      n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, 
      n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, 
      n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, 
      n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, 
      n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, 
      n2091, n2092, n2093, n2094, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
      n12, n13, n14, n15, n16, n17, n18, n19, n20, n2095, n2096, n2097, n2098, 
      n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, 
      n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, 
      n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, 
      n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, 
      n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, 
      n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, 
      n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, 
      n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, 
      n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, 
      n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, 
      n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, 
      n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, 
      n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, 
      n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, 
      n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, 
      n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, 
      n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, 
      n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, 
      n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, 
      n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, 
      n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, 
      n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, 
      n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, 
      n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, 
      n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, 
      n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, 
      n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, 
      n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, 
      n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, 
      n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, 
      n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, 
      n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, 
      n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, 
      n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, 
      n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, 
      n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, 
      n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, 
      n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, 
      n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, 
      n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, 
      n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, 
      n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, 
      n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, 
      n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, 
      n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, 
      n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, 
      n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, 
      n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, 
      n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, 
      n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, 
      n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, 
      n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, 
      n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, 
      n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, 
      n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, 
      n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, 
      n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, 
      n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, 
      n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, 
      n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, 
      n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, 
      n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, 
      n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, 
      n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, 
      n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, 
      n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, 
      n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, 
      n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, 
      n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, 
      n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, 
      n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, 
      n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, 
      n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, 
      n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, 
      n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, 
      n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, 
      n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, 
      n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, 
      n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, 
      n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, 
      n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, 
      n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, 
      n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, 
      n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, 
      n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, 
      n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, 
      n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, 
      n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, 
      n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, 
      n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, 
      n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, 
      n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, 
      n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, 
      n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, 
      n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, 
      n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, 
      n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, 
      n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, 
      n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, 
      n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, 
      n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, 
      n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, 
      n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, 
      n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, 
      n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, 
      n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, 
      n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, 
      n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, 
      n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, 
      n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, 
      n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, 
      n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, 
      n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, 
      n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, 
      n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, 
      n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, 
      n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, 
      n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, 
      n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, 
      n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, 
      n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, 
      n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, 
      n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, 
      n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, 
      n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, 
      n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, 
      n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, 
      n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, 
      n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, 
      n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, 
      n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, 
      n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, 
      n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, 
      n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, 
      n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, 
      n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, 
      n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, 
      n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, 
      n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, 
      n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, 
      n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, 
      n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, 
      n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, 
      n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, 
      n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, 
      n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, 
      n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, 
      n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, 
      n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, 
      n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, 
      n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, 
      n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, 
      n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, 
      n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, 
      n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, 
      n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, 
      n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, 
      n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, 
      n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, 
      n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, 
      n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, 
      n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, 
      n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, 
      n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, 
      n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, 
      n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, 
      n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, 
      n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, 
      n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, 
      n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, 
      n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, 
      n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, 
      n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, 
      n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, 
      n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, 
      n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, 
      n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, 
      n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, 
      n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, 
      n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, 
      n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, 
      n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, 
      n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, 
      n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, 
      n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, 
      n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, 
      n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, 
      n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, 
      n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, 
      n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, 
      n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, 
      n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, 
      n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, 
      n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, 
      n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, 
      n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, 
      n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, 
      n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, 
      n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, 
      n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, 
      n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, 
      n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, 
      n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, 
      n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, 
      n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, 
      n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, 
      n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, 
      n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, 
      n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, 
      n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, 
      n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, 
      n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, 
      n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, 
      n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, 
      n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, 
      n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, 
      n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, 
      n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, 
      n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, 
      n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, 
      n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, 
      n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, 
      n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, 
      n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, 
      n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, 
      n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, 
      n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, 
      n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, 
      n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, 
      n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, 
      n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, 
      n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, 
      n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, 
      n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, 
      n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, 
      n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, 
      n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, 
      n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, 
      n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, 
      n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, 
      n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, 
      n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, 
      n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, 
      n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, 
      n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, 
      n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, 
      n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, 
      n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, 
      n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, 
      n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, 
      n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, 
      n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, 
      n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, 
      n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, 
      n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, 
      n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, 
      n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, 
      n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, 
      n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, 
      n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, 
      n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, 
      n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, 
      n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, 
      n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, 
      n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, 
      n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, 
      n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, 
      n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, 
      n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, 
      n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, 
      n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, 
      n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, 
      n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, 
      n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, 
      n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, 
      n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, 
      n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, 
      n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, 
      n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, 
      n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, 
      n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, 
      n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, 
      n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, 
      n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, 
      n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, 
      n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, 
      n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, 
      n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, 
      n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, 
      n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, 
      n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, 
      n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, 
      n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, 
      n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, 
      n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, 
      n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, 
      n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, 
      n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, 
      n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, 
      n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, 
      n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, 
      n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, 
      n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, 
      n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, 
      n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, 
      n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, 
      n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, 
      n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, 
      n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, 
      n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, 
      n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, 
      n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, 
      n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, 
      n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, 
      n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, 
      n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, 
      n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, 
      n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, 
      n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, 
      n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, 
      n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, 
      n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, 
      n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, 
      n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, 
      n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, 
      n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, 
      n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, 
      n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, 
      n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, 
      n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, 
      n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, 
      n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, 
      n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, 
      n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, 
      n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, 
      n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, 
      n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, 
      n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, 
      n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, 
      n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, 
      n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, 
      n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, 
      n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, 
      n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, 
      n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, 
      n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, 
      n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, 
      n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, 
      n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, 
      n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, 
      n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, 
      n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n_1029, 
      n_1030, n_1031, n_1032, n_1033, n_1034, n_1035, n_1036, n_1037, n_1038, 
      n_1039, n_1040, n_1041, n_1042, n_1043, n_1044, n_1045, n_1046, n_1047, 
      n_1048, n_1049, n_1050, n_1051, n_1052, n_1053, n_1054, n_1055, n_1056, 
      n_1057, n_1058, n_1059, n_1060, n_1061, n_1062, n_1063, n_1064, n_1065, 
      n_1066, n_1067, n_1068, n_1069, n_1070, n_1071, n_1072, n_1073, n_1074, 
      n_1075, n_1076, n_1077, n_1078, n_1079, n_1080, n_1081, n_1082, n_1083, 
      n_1084, n_1085, n_1086, n_1087, n_1088, n_1089, n_1090, n_1091, n_1092, 
      n_1093, n_1094, n_1095, n_1096, n_1097, n_1098, n_1099, n_1100, n_1101, 
      n_1102, n_1103, n_1104, n_1105, n_1106, n_1107, n_1108, n_1109, n_1110, 
      n_1111, n_1112, n_1113, n_1114, n_1115, n_1116, n_1117, n_1118, n_1119, 
      n_1120, n_1121, n_1122, n_1123, n_1124, n_1125, n_1126, n_1127, n_1128, 
      n_1129, n_1130, n_1131, n_1132, n_1133, n_1134, n_1135, n_1136, n_1137, 
      n_1138, n_1139, n_1140, n_1141, n_1142, n_1143, n_1144, n_1145, n_1146, 
      n_1147, n_1148, n_1149, n_1150, n_1151, n_1152, n_1153, n_1154, n_1155, 
      n_1156, n_1157, n_1158, n_1159, n_1160, n_1161, n_1162, n_1163, n_1164, 
      n_1165, n_1166, n_1167, n_1168, n_1169, n_1170, n_1171, n_1172, n_1173, 
      n_1174, n_1175, n_1176, n_1177, n_1178, n_1179, n_1180, n_1181, n_1182, 
      n_1183, n_1184, n_1185, n_1186, n_1187, n_1188, n_1189, n_1190, n_1191, 
      n_1192, n_1193, n_1194, n_1195, n_1196, n_1197, n_1198, n_1199, n_1200, 
      n_1201, n_1202, n_1203, n_1204, n_1205, n_1206, n_1207, n_1208, n_1209, 
      n_1210, n_1211, n_1212, n_1213, n_1214, n_1215, n_1216, n_1217, n_1218, 
      n_1219, n_1220, n_1221, n_1222, n_1223, n_1224, n_1225, n_1226, n_1227, 
      n_1228, n_1229, n_1230, n_1231, n_1232, n_1233, n_1234, n_1235, n_1236, 
      n_1237, n_1238, n_1239, n_1240, n_1241, n_1242, n_1243, n_1244, n_1245, 
      n_1246, n_1247, n_1248, n_1249, n_1250, n_1251, n_1252, n_1253, n_1254, 
      n_1255, n_1256, n_1257, n_1258, n_1259, n_1260, n_1261, n_1262, n_1263, 
      n_1264, n_1265, n_1266, n_1267, n_1268, n_1269, n_1270, n_1271, n_1272, 
      n_1273, n_1274, n_1275, n_1276, n_1277, n_1278, n_1279, n_1280, n_1281, 
      n_1282, n_1283, n_1284, n_1285, n_1286, n_1287, n_1288, n_1289, n_1290, 
      n_1291, n_1292, n_1293, n_1294, n_1295, n_1296, n_1297, n_1298, n_1299, 
      n_1300, n_1301, n_1302, n_1303, n_1304, n_1305, n_1306, n_1307, n_1308, 
      n_1309, n_1310, n_1311, n_1312, n_1313, n_1314, n_1315, n_1316, n_1317, 
      n_1318, n_1319, n_1320, n_1321, n_1322, n_1323, n_1324, n_1325, n_1326, 
      n_1327, n_1328, n_1329, n_1330, n_1331, n_1332, n_1333, n_1334, n_1335, 
      n_1336, n_1337, n_1338, n_1339, n_1340, n_1341, n_1342, n_1343, n_1344, 
      n_1345, n_1346, n_1347, n_1348, n_1349, n_1350, n_1351, n_1352, n_1353, 
      n_1354, n_1355, n_1356, n_1357, n_1358, n_1359, n_1360, n_1361, n_1362, 
      n_1363, n_1364, n_1365, n_1366, n_1367, n_1368, n_1369, n_1370, n_1371, 
      n_1372, n_1373, n_1374, n_1375, n_1376, n_1377, n_1378, n_1379, n_1380, 
      n_1381, n_1382, n_1383, n_1384, n_1385, n_1386, n_1387, n_1388, n_1389, 
      n_1390, n_1391, n_1392, n_1393, n_1394, n_1395, n_1396, n_1397, n_1398, 
      n_1399, n_1400, n_1401, n_1402, n_1403, n_1404, n_1405, n_1406, n_1407, 
      n_1408, n_1409, n_1410, n_1411, n_1412, n_1413, n_1414, n_1415, n_1416, 
      n_1417, n_1418, n_1419, n_1420, n_1421, n_1422, n_1423, n_1424, n_1425, 
      n_1426, n_1427, n_1428, n_1429, n_1430, n_1431, n_1432, n_1433, n_1434, 
      n_1435, n_1436, n_1437, n_1438, n_1439, n_1440, n_1441, n_1442, n_1443, 
      n_1444, n_1445, n_1446, n_1447, n_1448, n_1449, n_1450, n_1451, n_1452, 
      n_1453, n_1454, n_1455, n_1456, n_1457, n_1458, n_1459, n_1460, n_1461, 
      n_1462, n_1463, n_1464, n_1465, n_1466, n_1467, n_1468, n_1469, n_1470, 
      n_1471, n_1472, n_1473, n_1474, n_1475, n_1476, n_1477, n_1478, n_1479, 
      n_1480, n_1481, n_1482, n_1483, n_1484, n_1485, n_1486, n_1487, n_1488, 
      n_1489, n_1490, n_1491, n_1492, n_1493, n_1494, n_1495, n_1496, n_1497, 
      n_1498, n_1499, n_1500, n_1501, n_1502, n_1503, n_1504, n_1505, n_1506, 
      n_1507, n_1508, n_1509, n_1510, n_1511, n_1512, n_1513, n_1514, n_1515, 
      n_1516, n_1517, n_1518, n_1519, n_1520, n_1521, n_1522, n_1523, n_1524, 
      n_1525, n_1526, n_1527, n_1528, n_1529, n_1530, n_1531, n_1532, n_1533, 
      n_1534, n_1535, n_1536, n_1537, n_1538, n_1539, n_1540, n_1541, n_1542, 
      n_1543, n_1544, n_1545, n_1546, n_1547, n_1548, n_1549, n_1550, n_1551, 
      n_1552, n_1553, n_1554, n_1555, n_1556, n_1557, n_1558, n_1559, n_1560, 
      n_1561, n_1562, n_1563, n_1564, n_1565, n_1566, n_1567, n_1568, n_1569, 
      n_1570, n_1571, n_1572, n_1573, n_1574, n_1575, n_1576, n_1577, n_1578, 
      n_1579, n_1580, n_1581, n_1582, n_1583, n_1584, n_1585, n_1586, n_1587, 
      n_1588, n_1589, n_1590, n_1591, n_1592, n_1593, n_1594, n_1595, n_1596, 
      n_1597, n_1598, n_1599, n_1600, n_1601, n_1602, n_1603, n_1604, n_1605, 
      n_1606, n_1607, n_1608, n_1609, n_1610, n_1611, n_1612, n_1613, n_1614, 
      n_1615, n_1616, n_1617, n_1618, n_1619, n_1620, n_1621, n_1622, n_1623, 
      n_1624, n_1625, n_1626, n_1627, n_1628, n_1629, n_1630, n_1631, n_1632, 
      n_1633, n_1634, n_1635, n_1636, n_1637, n_1638, n_1639, n_1640, n_1641, 
      n_1642, n_1643, n_1644, n_1645, n_1646, n_1647, n_1648, n_1649, n_1650, 
      n_1651, n_1652, n_1653, n_1654, n_1655, n_1656, n_1657, n_1658, n_1659, 
      n_1660, n_1661, n_1662, n_1663, n_1664, n_1665, n_1666, n_1667, n_1668, 
      n_1669, n_1670, n_1671, n_1672, n_1673, n_1674, n_1675, n_1676, n_1677, 
      n_1678, n_1679, n_1680, n_1681, n_1682, n_1683, n_1684, n_1685, n_1686, 
      n_1687, n_1688, n_1689, n_1690, n_1691, n_1692, n_1693, n_1694, n_1695, 
      n_1696, n_1697, n_1698, n_1699, n_1700, n_1701, n_1702, n_1703, n_1704, 
      n_1705, n_1706, n_1707, n_1708, n_1709, n_1710, n_1711, n_1712, n_1713, 
      n_1714, n_1715, n_1716, n_1717, n_1718, n_1719, n_1720, n_1721, n_1722, 
      n_1723, n_1724, n_1725, n_1726, n_1727, n_1728, n_1729, n_1730, n_1731, 
      n_1732, n_1733, n_1734, n_1735, n_1736, n_1737, n_1738, n_1739, n_1740, 
      n_1741, n_1742, n_1743, n_1744, n_1745, n_1746, n_1747, n_1748, n_1749, 
      n_1750, n_1751, n_1752, n_1753, n_1754, n_1755, n_1756, n_1757, n_1758, 
      n_1759, n_1760, n_1761, n_1762, n_1763, n_1764, n_1765, n_1766, n_1767, 
      n_1768, n_1769, n_1770, n_1771, n_1772, n_1773, n_1774, n_1775, n_1776, 
      n_1777, n_1778, n_1779, n_1780, n_1781, n_1782, n_1783, n_1784, n_1785, 
      n_1786, n_1787, n_1788, n_1789, n_1790, n_1791, n_1792, n_1793, n_1794, 
      n_1795, n_1796, n_1797, n_1798, n_1799, n_1800, n_1801, n_1802, n_1803, 
      n_1804, n_1805, n_1806, n_1807, n_1808, n_1809, n_1810, n_1811, n_1812, 
      n_1813, n_1814, n_1815, n_1816, n_1817, n_1818, n_1819, n_1820, n_1821, 
      n_1822, n_1823, n_1824, n_1825, n_1826, n_1827, n_1828, n_1829, n_1830, 
      n_1831, n_1832, n_1833, n_1834, n_1835, n_1836, n_1837, n_1838, n_1839, 
      n_1840, n_1841, n_1842, n_1843, n_1844, n_1845, n_1846, n_1847, n_1848, 
      n_1849, n_1850, n_1851, n_1852, n_1853, n_1854, n_1855, n_1856, n_1857, 
      n_1858, n_1859, n_1860, n_1861, n_1862, n_1863, n_1864, n_1865, n_1866, 
      n_1867, n_1868, n_1869, n_1870, n_1871, n_1872, n_1873, n_1874, n_1875, 
      n_1876, n_1877, n_1878, n_1879, n_1880, n_1881, n_1882, n_1883, n_1884, 
      n_1885, n_1886, n_1887, n_1888, n_1889, n_1890, n_1891, n_1892, n_1893, 
      n_1894, n_1895, n_1896, n_1897, n_1898, n_1899, n_1900, n_1901, n_1902, 
      n_1903, n_1904, n_1905, n_1906, n_1907, n_1908, n_1909, n_1910, n_1911, 
      n_1912, n_1913, n_1914, n_1915, n_1916, n_1917, n_1918, n_1919, n_1920, 
      n_1921, n_1922, n_1923, n_1924, n_1925, n_1926, n_1927, n_1928, n_1929, 
      n_1930, n_1931, n_1932, n_1933, n_1934, n_1935, n_1936, n_1937, n_1938, 
      n_1939, n_1940, n_1941, n_1942, n_1943, n_1944, n_1945, n_1946, n_1947, 
      n_1948, n_1949, n_1950, n_1951, n_1952, n_1953, n_1954, n_1955, n_1956, 
      n_1957, n_1958, n_1959, n_1960, n_1961, n_1962, n_1963, n_1964, n_1965, 
      n_1966, n_1967, n_1968, n_1969, n_1970, n_1971, n_1972, n_1973, n_1974, 
      n_1975, n_1976, n_1977, n_1978, n_1979, n_1980, n_1981, n_1982, n_1983, 
      n_1984, n_1985, n_1986, n_1987, n_1988, n_1989, n_1990, n_1991, n_1992, 
      n_1993, n_1994, n_1995, n_1996, n_1997, n_1998, n_1999, n_2000, n_2001, 
      n_2002, n_2003, n_2004, n_2005, n_2006, n_2007, n_2008, n_2009, n_2010, 
      n_2011, n_2012, n_2013, n_2014, n_2015, n_2016, n_2017, n_2018, n_2019, 
      n_2020, n_2021, n_2022, n_2023, n_2024, n_2025, n_2026, n_2027, n_2028, 
      n_2029, n_2030, n_2031, n_2032, n_2033, n_2034, n_2035, n_2036, n_2037, 
      n_2038, n_2039, n_2040, n_2041, n_2042, n_2043, n_2044, n_2045, n_2046, 
      n_2047, n_2048, n_2049, n_2050, n_2051, n_2052, n_2053, n_2054, n_2055, 
      n_2056, n_2057, n_2058, n_2059, n_2060, n_2061, n_2062, n_2063, n_2064, 
      n_2065, n_2066, n_2067, n_2068, n_2069, n_2070, n_2071, n_2072, n_2073, 
      n_2074, n_2075, n_2076, n_2077, n_2078, n_2079, n_2080, n_2081, n_2082, 
      n_2083, n_2084, n_2085, n_2086, n_2087, n_2088, n_2089, n_2090, n_2091, 
      n_2092, n_2093, n_2094, n_2095, n_2096, n_2097, n_2098, n_2099, n_2100, 
      n_2101, n_2102, n_2103, n_2104, n_2105, n_2106, n_2107, n_2108, n_2109, 
      n_2110, n_2111, n_2112, n_2113, n_2114, n_2115, n_2116, n_2117, n_2118, 
      n_2119, n_2120, n_2121, n_2122, n_2123, n_2124, n_2125, n_2126, n_2127, 
      n_2128, n_2129, n_2130, n_2131, n_2132, n_2133, n_2134, n_2135, n_2136, 
      n_2137, n_2138, n_2139, n_2140, n_2141, n_2142, n_2143, n_2144, n_2145, 
      n_2146, n_2147, n_2148, n_2149, n_2150, n_2151, n_2152, n_2153, n_2154, 
      n_2155, n_2156, n_2157, n_2158, n_2159, n_2160, n_2161, n_2162, n_2163, 
      n_2164, n_2165, n_2166, n_2167, n_2168, n_2169, n_2170, n_2171, n_2172, 
      n_2173, n_2174, n_2175, n_2176, n_2177, n_2178, n_2179, n_2180, n_2181, 
      n_2182, n_2183, n_2184, n_2185, n_2186, n_2187, n_2188, n_2189, n_2190, 
      n_2191, n_2192, n_2193, n_2194, n_2195, n_2196, n_2197, n_2198, n_2199, 
      n_2200, n_2201, n_2202, n_2203, n_2204, n_2205, n_2206, n_2207, n_2208, 
      n_2209, n_2210, n_2211, n_2212, n_2213, n_2214, n_2215, n_2216, n_2217, 
      n_2218, n_2219, n_2220, n_2221, n_2222, n_2223, n_2224, n_2225, n_2226, 
      n_2227, n_2228, n_2229, n_2230, n_2231, n_2232, n_2233, n_2234, n_2235, 
      n_2236, n_2237, n_2238, n_2239, n_2240, n_2241, n_2242, n_2243, n_2244, 
      n_2245, n_2246, n_2247, n_2248, n_2249, n_2250, n_2251, n_2252, n_2253, 
      n_2254, n_2255, n_2256, n_2257, n_2258, n_2259, n_2260, n_2261, n_2262, 
      n_2263, n_2264, n_2265, n_2266, n_2267, n_2268, n_2269, n_2270, n_2271, 
      n_2272, n_2273, n_2274, n_2275, n_2276, n_2277, n_2278, n_2279, n_2280, 
      n_2281, n_2282, n_2283, n_2284, n_2285, n_2286, n_2287, n_2288, n_2289, 
      n_2290, n_2291, n_2292, n_2293, n_2294, n_2295, n_2296, n_2297, n_2298, 
      n_2299, n_2300, n_2301, n_2302, n_2303, n_2304, n_2305, n_2306, n_2307, 
      n_2308, n_2309, n_2310, n_2311, n_2312, n_2313, n_2314, n_2315, n_2316, 
      n_2317, n_2318, n_2319, n_2320, n_2321, n_2322, n_2323, n_2324, n_2325, 
      n_2326, n_2327, n_2328, n_2329, n_2330, n_2331, n_2332, n_2333, n_2334, 
      n_2335, n_2336, n_2337, n_2338, n_2339, n_2340, n_2341, n_2342, n_2343, 
      n_2344, n_2345, n_2346, n_2347, n_2348, n_2349, n_2350, n_2351, n_2352, 
      n_2353, n_2354, n_2355, n_2356, n_2357, n_2358, n_2359, n_2360, n_2361, 
      n_2362, n_2363, n_2364, n_2365, n_2366, n_2367, n_2368, n_2369, n_2370, 
      n_2371, n_2372, n_2373, n_2374, n_2375, n_2376, n_2377, n_2378, n_2379, 
      n_2380, n_2381, n_2382, n_2383, n_2384, n_2385, n_2386, n_2387, n_2388, 
      n_2389, n_2390, n_2391, n_2392, n_2393, n_2394, n_2395, n_2396, n_2397, 
      n_2398, n_2399, n_2400, n_2401, n_2402, n_2403, n_2404, n_2405, n_2406, 
      n_2407, n_2408, n_2409, n_2410, n_2411, n_2412, n_2413, n_2414, n_2415, 
      n_2416, n_2417, n_2418, n_2419, n_2420, n_2421, n_2422, n_2423, n_2424, 
      n_2425, n_2426, n_2427, n_2428, n_2429, n_2430, n_2431, n_2432, n_2433, 
      n_2434, n_2435, n_2436, n_2437, n_2438, n_2439, n_2440, n_2441, n_2442, 
      n_2443, n_2444, n_2445, n_2446, n_2447, n_2448, n_2449, n_2450, n_2451, 
      n_2452, n_2453, n_2454, n_2455, n_2456, n_2457, n_2458, n_2459, n_2460, 
      n_2461, n_2462, n_2463, n_2464, n_2465, n_2466, n_2467, n_2468, n_2469, 
      n_2470, n_2471, n_2472, n_2473, n_2474, n_2475, n_2476, n_2477, n_2478, 
      n_2479, n_2480, n_2481, n_2482, n_2483, n_2484, n_2485, n_2486, n_2487, 
      n_2488, n_2489, n_2490, n_2491, n_2492, n_2493, n_2494, n_2495, n_2496, 
      n_2497, n_2498, n_2499, n_2500, n_2501, n_2502, n_2503, n_2504, n_2505, 
      n_2506, n_2507, n_2508, n_2509, n_2510, n_2511, n_2512, n_2513, n_2514, 
      n_2515, n_2516, n_2517, n_2518, n_2519, n_2520, n_2521, n_2522, n_2523, 
      n_2524, n_2525, n_2526, n_2527, n_2528, n_2529, n_2530, n_2531, n_2532, 
      n_2533, n_2534, n_2535, n_2536, n_2537, n_2538, n_2539, n_2540, n_2541, 
      n_2542, n_2543, n_2544, n_2545, n_2546, n_2547, n_2548, n_2549, n_2550, 
      n_2551, n_2552, n_2553, n_2554, n_2555, n_2556, n_2557, n_2558, n_2559, 
      n_2560, n_2561, n_2562, n_2563, n_2564, n_2565, n_2566, n_2567, n_2568, 
      n_2569, n_2570, n_2571, n_2572, n_2573, n_2574, n_2575, n_2576, n_2577, 
      n_2578, n_2579, n_2580, n_2581, n_2582, n_2583, n_2584, n_2585, n_2586, 
      n_2587, n_2588, n_2589, n_2590, n_2591, n_2592, n_2593, n_2594, n_2595, 
      n_2596, n_2597, n_2598, n_2599, n_2600, n_2601, n_2602, n_2603, n_2604, 
      n_2605, n_2606, n_2607, n_2608, n_2609, n_2610, n_2611, n_2612, n_2613, 
      n_2614, n_2615, n_2616, n_2617, n_2618, n_2619, n_2620, n_2621, n_2622, 
      n_2623, n_2624, n_2625, n_2626, n_2627, n_2628, n_2629, n_2630, n_2631, 
      n_2632, n_2633, n_2634, n_2635, n_2636, n_2637, n_2638, n_2639, n_2640, 
      n_2641, n_2642, n_2643, n_2644, n_2645, n_2646, n_2647, n_2648, n_2649, 
      n_2650, n_2651, n_2652, n_2653, n_2654, n_2655, n_2656, n_2657, n_2658, 
      n_2659, n_2660, n_2661, n_2662, n_2663, n_2664, n_2665, n_2666, n_2667, 
      n_2668, n_2669, n_2670, n_2671, n_2672, n_2673, n_2674, n_2675, n_2676, 
      n_2677, n_2678, n_2679, n_2680, n_2681, n_2682, n_2683, n_2684, n_2685, 
      n_2686, n_2687, n_2688, n_2689, n_2690, n_2691, n_2692, n_2693, n_2694, 
      n_2695, n_2696, n_2697, n_2698, n_2699, n_2700, n_2701, n_2702, n_2703, 
      n_2704, n_2705, n_2706, n_2707, n_2708, n_2709, n_2710, n_2711, n_2712, 
      n_2713, n_2714, n_2715, n_2716, n_2717, n_2718, n_2719, n_2720, n_2721, 
      n_2722, n_2723, n_2724, n_2725, n_2726, n_2727, n_2728, n_2729, n_2730, 
      n_2731, n_2732, n_2733, n_2734, n_2735, n_2736, n_2737, n_2738, n_2739, 
      n_2740, n_2741, n_2742, n_2743, n_2744, n_2745, n_2746, n_2747, n_2748, 
      n_2749, n_2750, n_2751, n_2752, n_2753, n_2754, n_2755, n_2756, n_2757, 
      n_2758, n_2759, n_2760, n_2761, n_2762, n_2763, n_2764, n_2765, n_2766, 
      n_2767, n_2768, n_2769, n_2770, n_2771, n_2772, n_2773, n_2774, n_2775, 
      n_2776, n_2777, n_2778, n_2779, n_2780, n_2781, n_2782, n_2783, n_2784, 
      n_2785, n_2786, n_2787, n_2788, n_2789, n_2790, n_2791, n_2792, n_2793, 
      n_2794, n_2795, n_2796, n_2797, n_2798, n_2799, n_2800, n_2801, n_2802, 
      n_2803, n_2804, n_2805, n_2806, n_2807, n_2808, n_2809, n_2810, n_2811, 
      n_2812, n_2813, n_2814, n_2815, n_2816, n_2817, n_2818, n_2819, n_2820, 
      n_2821, n_2822, n_2823, n_2824, n_2825, n_2826, n_2827, n_2828, n_2829, 
      n_2830, n_2831, n_2832, n_2833, n_2834, n_2835, n_2836, n_2837, n_2838, 
      n_2839, n_2840, n_2841, n_2842, n_2843, n_2844, n_2845, n_2846, n_2847, 
      n_2848, n_2849, n_2850, n_2851, n_2852, n_2853, n_2854, n_2855, n_2856, 
      n_2857, n_2858, n_2859, n_2860, n_2861, n_2862, n_2863, n_2864, n_2865, 
      n_2866, n_2867, n_2868, n_2869, n_2870, n_2871, n_2872, n_2873, n_2874, 
      n_2875, n_2876, n_2877, n_2878, n_2879, n_2880, n_2881, n_2882, n_2883, 
      n_2884, n_2885, n_2886, n_2887, n_2888, n_2889, n_2890, n_2891, n_2892, 
      n_2893, n_2894, n_2895, n_2896, n_2897, n_2898, n_2899, n_2900, n_2901, 
      n_2902, n_2903, n_2904, n_2905, n_2906, n_2907, n_2908, n_2909, n_2910, 
      n_2911, n_2912, n_2913, n_2914, n_2915, n_2916, n_2917, n_2918, n_2919, 
      n_2920, n_2921, n_2922, n_2923, n_2924, n_2925, n_2926, n_2927, n_2928, 
      n_2929, n_2930, n_2931, n_2932, n_2933, n_2934, n_2935, n_2936, n_2937, 
      n_2938, n_2939, n_2940, n_2941, n_2942, n_2943, n_2944, n_2945, n_2946, 
      n_2947, n_2948, n_2949, n_2950, n_2951, n_2952, n_2953, n_2954, n_2955, 
      n_2956, n_2957, n_2958, n_2959, n_2960, n_2961, n_2962, n_2963, n_2964, 
      n_2965, n_2966, n_2967, n_2968, n_2969, n_2970, n_2971, n_2972, n_2973, 
      n_2974, n_2975, n_2976, n_2977, n_2978, n_2979, n_2980, n_2981, n_2982, 
      n_2983, n_2984, n_2985, n_2986, n_2987, n_2988, n_2989, n_2990, n_2991, 
      n_2992, n_2993, n_2994, n_2995, n_2996, n_2997, n_2998, n_2999, n_3000, 
      n_3001, n_3002, n_3003, n_3004, n_3005, n_3006, n_3007, n_3008, n_3009, 
      n_3010, n_3011, n_3012, n_3013, n_3014, n_3015, n_3016, n_3017, n_3018, 
      n_3019, n_3020, n_3021, n_3022, n_3023, n_3024, n_3025, n_3026, n_3027, 
      n_3028, n_3029, n_3030, n_3031, n_3032, n_3033, n_3034, n_3035, n_3036, 
      n_3037, n_3038, n_3039, n_3040, n_3041, n_3042, n_3043, n_3044, n_3045, 
      n_3046, n_3047, n_3048, n_3049, n_3050, n_3051, n_3052, n_3053, n_3054, 
      n_3055, n_3056, n_3057, n_3058, n_3059, n_3060, n_3061, n_3062, n_3063, 
      n_3064, n_3065, n_3066, n_3067, n_3068, n_3069, n_3070, n_3071, n_3072, 
      n_3073, n_3074, n_3075, n_3076 : std_logic;

begin
   
   RAM_reg_0_127_inst : DFFX1 port map( D => n2094, CLK => n4781, Q => 
                           RAM_0_127_port, QN => n_1029);
   RAM_reg_0_126_inst : DFFX1 port map( D => n2093, CLK => n4781, Q => 
                           RAM_0_126_port, QN => n_1030);
   RAM_reg_0_125_inst : DFFX1 port map( D => n2092, CLK => n4781, Q => 
                           RAM_0_125_port, QN => n_1031);
   RAM_reg_0_124_inst : DFFX1 port map( D => n2091, CLK => n4781, Q => 
                           RAM_0_124_port, QN => n_1032);
   RAM_reg_0_123_inst : DFFX1 port map( D => n2090, CLK => n4781, Q => 
                           RAM_0_123_port, QN => n_1033);
   RAM_reg_0_122_inst : DFFX1 port map( D => n2089, CLK => n4781, Q => 
                           RAM_0_122_port, QN => n_1034);
   RAM_reg_0_121_inst : DFFX1 port map( D => n2088, CLK => n4781, Q => 
                           RAM_0_121_port, QN => n_1035);
   RAM_reg_0_120_inst : DFFX1 port map( D => n2087, CLK => n4781, Q => 
                           RAM_0_120_port, QN => n_1036);
   RAM_reg_0_119_inst : DFFX1 port map( D => n2086, CLK => n4781, Q => 
                           RAM_0_119_port, QN => n_1037);
   RAM_reg_0_118_inst : DFFX1 port map( D => n2085, CLK => n4781, Q => 
                           RAM_0_118_port, QN => n_1038);
   RAM_reg_0_117_inst : DFFX1 port map( D => n2084, CLK => n4781, Q => 
                           RAM_0_117_port, QN => n_1039);
   RAM_reg_0_116_inst : DFFX1 port map( D => n2083, CLK => n4781, Q => 
                           RAM_0_116_port, QN => n_1040);
   RAM_reg_0_115_inst : DFFX1 port map( D => n2082, CLK => n4782, Q => 
                           RAM_0_115_port, QN => n_1041);
   RAM_reg_0_114_inst : DFFX1 port map( D => n2081, CLK => n4782, Q => 
                           RAM_0_114_port, QN => n_1042);
   RAM_reg_0_113_inst : DFFX1 port map( D => n2080, CLK => n4782, Q => 
                           RAM_0_113_port, QN => n_1043);
   RAM_reg_0_112_inst : DFFX1 port map( D => n2079, CLK => n4782, Q => 
                           RAM_0_112_port, QN => n_1044);
   RAM_reg_0_111_inst : DFFX1 port map( D => n2078, CLK => n4782, Q => 
                           RAM_0_111_port, QN => n_1045);
   RAM_reg_0_110_inst : DFFX1 port map( D => n2077, CLK => n4782, Q => 
                           RAM_0_110_port, QN => n_1046);
   RAM_reg_0_109_inst : DFFX1 port map( D => n2076, CLK => n4782, Q => 
                           RAM_0_109_port, QN => n_1047);
   RAM_reg_0_108_inst : DFFX1 port map( D => n2075, CLK => n4782, Q => 
                           RAM_0_108_port, QN => n_1048);
   RAM_reg_0_107_inst : DFFX1 port map( D => n2074, CLK => n4782, Q => 
                           RAM_0_107_port, QN => n_1049);
   RAM_reg_0_106_inst : DFFX1 port map( D => n2073, CLK => n4782, Q => 
                           RAM_0_106_port, QN => n_1050);
   RAM_reg_0_105_inst : DFFX1 port map( D => n2072, CLK => n4782, Q => 
                           RAM_0_105_port, QN => n_1051);
   RAM_reg_0_104_inst : DFFX1 port map( D => n2071, CLK => n4782, Q => 
                           RAM_0_104_port, QN => n_1052);
   RAM_reg_0_103_inst : DFFX1 port map( D => n2070, CLK => n4783, Q => 
                           RAM_0_103_port, QN => n_1053);
   RAM_reg_0_102_inst : DFFX1 port map( D => n2069, CLK => n4783, Q => 
                           RAM_0_102_port, QN => n_1054);
   RAM_reg_0_101_inst : DFFX1 port map( D => n2068, CLK => n4783, Q => 
                           RAM_0_101_port, QN => n_1055);
   RAM_reg_0_100_inst : DFFX1 port map( D => n2067, CLK => n4783, Q => 
                           RAM_0_100_port, QN => n_1056);
   RAM_reg_0_99_inst : DFFX1 port map( D => n2066, CLK => n4783, Q => 
                           RAM_0_99_port, QN => n_1057);
   RAM_reg_0_98_inst : DFFX1 port map( D => n2065, CLK => n4783, Q => 
                           RAM_0_98_port, QN => n_1058);
   RAM_reg_0_97_inst : DFFX1 port map( D => n2064, CLK => n4783, Q => 
                           RAM_0_97_port, QN => n_1059);
   RAM_reg_0_96_inst : DFFX1 port map( D => n2063, CLK => n4783, Q => 
                           RAM_0_96_port, QN => n_1060);
   RAM_reg_0_95_inst : DFFX1 port map( D => n2062, CLK => n4778, Q => 
                           RAM_0_95_port, QN => n_1061);
   RAM_reg_0_94_inst : DFFX1 port map( D => n2061, CLK => n4778, Q => 
                           RAM_0_94_port, QN => n_1062);
   RAM_reg_0_93_inst : DFFX1 port map( D => n2060, CLK => n4778, Q => 
                           RAM_0_93_port, QN => n_1063);
   RAM_reg_0_92_inst : DFFX1 port map( D => n2059, CLK => n4778, Q => 
                           RAM_0_92_port, QN => n_1064);
   RAM_reg_0_91_inst : DFFX1 port map( D => n2058, CLK => n4778, Q => 
                           RAM_0_91_port, QN => n_1065);
   RAM_reg_0_90_inst : DFFX1 port map( D => n2057, CLK => n4778, Q => 
                           RAM_0_90_port, QN => n_1066);
   RAM_reg_0_89_inst : DFFX1 port map( D => n2056, CLK => n4778, Q => 
                           RAM_0_89_port, QN => n_1067);
   RAM_reg_0_88_inst : DFFX1 port map( D => n2055, CLK => n4778, Q => 
                           RAM_0_88_port, QN => n_1068);
   RAM_reg_0_87_inst : DFFX1 port map( D => n2054, CLK => n4778, Q => 
                           RAM_0_87_port, QN => n_1069);
   RAM_reg_0_86_inst : DFFX1 port map( D => n2053, CLK => n4778, Q => 
                           RAM_0_86_port, QN => n_1070);
   RAM_reg_0_85_inst : DFFX1 port map( D => n2052, CLK => n4778, Q => 
                           RAM_0_85_port, QN => n_1071);
   RAM_reg_0_84_inst : DFFX1 port map( D => n2051, CLK => n4778, Q => 
                           RAM_0_84_port, QN => n_1072);
   RAM_reg_0_83_inst : DFFX1 port map( D => n2050, CLK => n4779, Q => 
                           RAM_0_83_port, QN => n_1073);
   RAM_reg_0_82_inst : DFFX1 port map( D => n2049, CLK => n4779, Q => 
                           RAM_0_82_port, QN => n_1074);
   RAM_reg_0_81_inst : DFFX1 port map( D => n2048, CLK => n4779, Q => 
                           RAM_0_81_port, QN => n_1075);
   RAM_reg_0_80_inst : DFFX1 port map( D => n2047, CLK => n4779, Q => 
                           RAM_0_80_port, QN => n_1076);
   RAM_reg_0_79_inst : DFFX1 port map( D => n2046, CLK => n4779, Q => 
                           RAM_0_79_port, QN => n_1077);
   RAM_reg_0_78_inst : DFFX1 port map( D => n2045, CLK => n4779, Q => 
                           RAM_0_78_port, QN => n_1078);
   RAM_reg_0_77_inst : DFFX1 port map( D => n2044, CLK => n4779, Q => 
                           RAM_0_77_port, QN => n_1079);
   RAM_reg_0_76_inst : DFFX1 port map( D => n2043, CLK => n4779, Q => 
                           RAM_0_76_port, QN => n_1080);
   RAM_reg_0_75_inst : DFFX1 port map( D => n2042, CLK => n4779, Q => 
                           RAM_0_75_port, QN => n_1081);
   RAM_reg_0_74_inst : DFFX1 port map( D => n2041, CLK => n4779, Q => 
                           RAM_0_74_port, QN => n_1082);
   RAM_reg_0_73_inst : DFFX1 port map( D => n2040, CLK => n4779, Q => 
                           RAM_0_73_port, QN => n_1083);
   RAM_reg_0_72_inst : DFFX1 port map( D => n2039, CLK => n4779, Q => 
                           RAM_0_72_port, QN => n_1084);
   RAM_reg_0_71_inst : DFFX1 port map( D => n2038, CLK => n4780, Q => 
                           RAM_0_71_port, QN => n_1085);
   RAM_reg_0_70_inst : DFFX1 port map( D => n2037, CLK => n4780, Q => 
                           RAM_0_70_port, QN => n_1086);
   RAM_reg_0_69_inst : DFFX1 port map( D => n2036, CLK => n4780, Q => 
                           RAM_0_69_port, QN => n_1087);
   RAM_reg_0_68_inst : DFFX1 port map( D => n2035, CLK => n4780, Q => 
                           RAM_0_68_port, QN => n_1088);
   RAM_reg_0_67_inst : DFFX1 port map( D => n2034, CLK => n4780, Q => 
                           RAM_0_67_port, QN => n_1089);
   RAM_reg_0_66_inst : DFFX1 port map( D => n2033, CLK => n4780, Q => 
                           RAM_0_66_port, QN => n_1090);
   RAM_reg_0_65_inst : DFFX1 port map( D => n2032, CLK => n4780, Q => 
                           RAM_0_65_port, QN => n_1091);
   RAM_reg_0_64_inst : DFFX1 port map( D => n2031, CLK => n4780, Q => 
                           RAM_0_64_port, QN => n_1092);
   RAM_reg_0_63_inst : DFFX1 port map( D => n2030, CLK => n4780, Q => 
                           RAM_0_63_port, QN => n_1093);
   RAM_reg_0_62_inst : DFFX1 port map( D => n2029, CLK => n4780, Q => 
                           RAM_0_62_port, QN => n_1094);
   RAM_reg_0_61_inst : DFFX1 port map( D => n2028, CLK => n4780, Q => 
                           RAM_0_61_port, QN => n_1095);
   RAM_reg_0_60_inst : DFFX1 port map( D => n2027, CLK => n4780, Q => 
                           RAM_0_60_port, QN => n_1096);
   RAM_reg_0_59_inst : DFFX1 port map( D => n2026, CLK => n4775, Q => 
                           RAM_0_59_port, QN => n_1097);
   RAM_reg_0_58_inst : DFFX1 port map( D => n2025, CLK => n4775, Q => 
                           RAM_0_58_port, QN => n_1098);
   RAM_reg_0_57_inst : DFFX1 port map( D => n2024, CLK => n4775, Q => 
                           RAM_0_57_port, QN => n_1099);
   RAM_reg_0_56_inst : DFFX1 port map( D => n2023, CLK => n4775, Q => 
                           RAM_0_56_port, QN => n_1100);
   RAM_reg_0_55_inst : DFFX1 port map( D => n2022, CLK => n4775, Q => 
                           RAM_0_55_port, QN => n_1101);
   RAM_reg_0_54_inst : DFFX1 port map( D => n2021, CLK => n4775, Q => 
                           RAM_0_54_port, QN => n_1102);
   RAM_reg_0_53_inst : DFFX1 port map( D => n2020, CLK => n4775, Q => 
                           RAM_0_53_port, QN => n_1103);
   RAM_reg_0_52_inst : DFFX1 port map( D => n2019, CLK => n4775, Q => 
                           RAM_0_52_port, QN => n_1104);
   RAM_reg_0_51_inst : DFFX1 port map( D => n2018, CLK => n4775, Q => 
                           RAM_0_51_port, QN => n_1105);
   RAM_reg_0_50_inst : DFFX1 port map( D => n2017, CLK => n4775, Q => 
                           RAM_0_50_port, QN => n_1106);
   RAM_reg_0_49_inst : DFFX1 port map( D => n2016, CLK => n4775, Q => 
                           RAM_0_49_port, QN => n_1107);
   RAM_reg_0_48_inst : DFFX1 port map( D => n2015, CLK => n4775, Q => 
                           RAM_0_48_port, QN => n_1108);
   RAM_reg_0_47_inst : DFFX1 port map( D => n2014, CLK => n4776, Q => 
                           RAM_0_47_port, QN => n_1109);
   RAM_reg_0_46_inst : DFFX1 port map( D => n2013, CLK => n4776, Q => 
                           RAM_0_46_port, QN => n_1110);
   RAM_reg_0_45_inst : DFFX1 port map( D => n2012, CLK => n4776, Q => 
                           RAM_0_45_port, QN => n_1111);
   RAM_reg_0_44_inst : DFFX1 port map( D => n2011, CLK => n4776, Q => 
                           RAM_0_44_port, QN => n_1112);
   RAM_reg_0_43_inst : DFFX1 port map( D => n2010, CLK => n4776, Q => 
                           RAM_0_43_port, QN => n_1113);
   RAM_reg_0_42_inst : DFFX1 port map( D => n2009, CLK => n4776, Q => 
                           RAM_0_42_port, QN => n_1114);
   RAM_reg_0_41_inst : DFFX1 port map( D => n2008, CLK => n4776, Q => 
                           RAM_0_41_port, QN => n_1115);
   RAM_reg_0_40_inst : DFFX1 port map( D => n2007, CLK => n4776, Q => 
                           RAM_0_40_port, QN => n_1116);
   RAM_reg_0_39_inst : DFFX1 port map( D => n2006, CLK => n4776, Q => 
                           RAM_0_39_port, QN => n_1117);
   RAM_reg_0_38_inst : DFFX1 port map( D => n2005, CLK => n4776, Q => 
                           RAM_0_38_port, QN => n_1118);
   RAM_reg_0_37_inst : DFFX1 port map( D => n2004, CLK => n4776, Q => 
                           RAM_0_37_port, QN => n_1119);
   RAM_reg_0_36_inst : DFFX1 port map( D => n2003, CLK => n4776, Q => 
                           RAM_0_36_port, QN => n_1120);
   RAM_reg_0_35_inst : DFFX1 port map( D => n2002, CLK => n4777, Q => 
                           RAM_0_35_port, QN => n_1121);
   RAM_reg_0_34_inst : DFFX1 port map( D => n2001, CLK => n4777, Q => 
                           RAM_0_34_port, QN => n_1122);
   RAM_reg_0_33_inst : DFFX1 port map( D => n2000, CLK => n4777, Q => 
                           RAM_0_33_port, QN => n_1123);
   RAM_reg_0_32_inst : DFFX1 port map( D => n1999, CLK => n4777, Q => 
                           RAM_0_32_port, QN => n_1124);
   RAM_reg_0_31_inst : DFFX1 port map( D => n1998, CLK => n4777, Q => 
                           RAM_0_31_port, QN => n_1125);
   RAM_reg_0_30_inst : DFFX1 port map( D => n1997, CLK => n4777, Q => 
                           RAM_0_30_port, QN => n_1126);
   RAM_reg_0_29_inst : DFFX1 port map( D => n1996, CLK => n4777, Q => 
                           RAM_0_29_port, QN => n_1127);
   RAM_reg_0_28_inst : DFFX1 port map( D => n1995, CLK => n4777, Q => 
                           RAM_0_28_port, QN => n_1128);
   RAM_reg_0_27_inst : DFFX1 port map( D => n1994, CLK => n4777, Q => 
                           RAM_0_27_port, QN => n_1129);
   RAM_reg_0_26_inst : DFFX1 port map( D => n1993, CLK => n4777, Q => 
                           RAM_0_26_port, QN => n_1130);
   RAM_reg_0_25_inst : DFFX1 port map( D => n1992, CLK => n4777, Q => 
                           RAM_0_25_port, QN => n_1131);
   RAM_reg_0_24_inst : DFFX1 port map( D => n1991, CLK => n4777, Q => 
                           RAM_0_24_port, QN => n_1132);
   RAM_reg_0_23_inst : DFFX1 port map( D => n1990, CLK => n4789, Q => 
                           RAM_0_23_port, QN => n_1133);
   RAM_reg_0_22_inst : DFFX1 port map( D => n1989, CLK => n4789, Q => 
                           RAM_0_22_port, QN => n_1134);
   RAM_reg_0_21_inst : DFFX1 port map( D => n1988, CLK => n4789, Q => 
                           RAM_0_21_port, QN => n_1135);
   RAM_reg_0_20_inst : DFFX1 port map( D => n1987, CLK => n4789, Q => 
                           RAM_0_20_port, QN => n_1136);
   RAM_reg_0_19_inst : DFFX1 port map( D => n1986, CLK => n4790, Q => 
                           RAM_0_19_port, QN => n_1137);
   RAM_reg_0_18_inst : DFFX1 port map( D => n1985, CLK => n4790, Q => 
                           RAM_0_18_port, QN => n_1138);
   RAM_reg_0_17_inst : DFFX1 port map( D => n1984, CLK => n4790, Q => 
                           RAM_0_17_port, QN => n_1139);
   RAM_reg_0_16_inst : DFFX1 port map( D => n1983, CLK => n4790, Q => 
                           RAM_0_16_port, QN => n_1140);
   RAM_reg_0_15_inst : DFFX1 port map( D => n1982, CLK => n4790, Q => 
                           RAM_0_15_port, QN => n_1141);
   RAM_reg_0_14_inst : DFFX1 port map( D => n1981, CLK => n4790, Q => 
                           RAM_0_14_port, QN => n_1142);
   RAM_reg_0_13_inst : DFFX1 port map( D => n1980, CLK => n4790, Q => 
                           RAM_0_13_port, QN => n_1143);
   RAM_reg_0_12_inst : DFFX1 port map( D => n1979, CLK => n4790, Q => 
                           RAM_0_12_port, QN => n_1144);
   RAM_reg_0_11_inst : DFFX1 port map( D => n1978, CLK => n4790, Q => 
                           RAM_0_11_port, QN => n_1145);
   RAM_reg_0_10_inst : DFFX1 port map( D => n1977, CLK => n4790, Q => 
                           RAM_0_10_port, QN => n_1146);
   RAM_reg_0_9_inst : DFFX1 port map( D => n1976, CLK => n4790, Q => 
                           RAM_0_9_port, QN => n_1147);
   RAM_reg_0_8_inst : DFFX1 port map( D => n1975, CLK => n4790, Q => 
                           RAM_0_8_port, QN => n_1148);
   RAM_reg_0_7_inst : DFFX1 port map( D => n1974, CLK => n4791, Q => 
                           RAM_0_7_port, QN => n_1149);
   RAM_reg_0_6_inst : DFFX1 port map( D => n1973, CLK => n4791, Q => 
                           RAM_0_6_port, QN => n_1150);
   RAM_reg_0_5_inst : DFFX1 port map( D => n1972, CLK => n4791, Q => 
                           RAM_0_5_port, QN => n_1151);
   RAM_reg_0_4_inst : DFFX1 port map( D => n1971, CLK => n4791, Q => 
                           RAM_0_4_port, QN => n_1152);
   RAM_reg_0_3_inst : DFFX1 port map( D => n1970, CLK => n4791, Q => 
                           RAM_0_3_port, QN => n_1153);
   RAM_reg_0_2_inst : DFFX1 port map( D => n1969, CLK => n4791, Q => 
                           RAM_0_2_port, QN => n_1154);
   RAM_reg_0_1_inst : DFFX1 port map( D => n1968, CLK => n4791, Q => 
                           RAM_0_1_port, QN => n_1155);
   RAM_reg_0_0_inst : DFFX1 port map( D => n1967, CLK => n4791, Q => 
                           RAM_0_0_port, QN => n_1156);
   RAM_reg_1_127_inst : DFFX1 port map( D => n1966, CLK => n4791, Q => 
                           RAM_1_127_port, QN => n_1157);
   RAM_reg_1_126_inst : DFFX1 port map( D => n1965, CLK => n4791, Q => 
                           RAM_1_126_port, QN => n_1158);
   RAM_reg_1_125_inst : DFFX1 port map( D => n1964, CLK => n4791, Q => 
                           RAM_1_125_port, QN => n_1159);
   RAM_reg_1_124_inst : DFFX1 port map( D => n1963, CLK => n4791, Q => 
                           RAM_1_124_port, QN => n_1160);
   RAM_reg_1_123_inst : DFFX1 port map( D => n1962, CLK => n4792, Q => 
                           RAM_1_123_port, QN => n_1161);
   RAM_reg_1_122_inst : DFFX1 port map( D => n1961, CLK => n4792, Q => 
                           RAM_1_122_port, QN => n_1162);
   RAM_reg_1_121_inst : DFFX1 port map( D => n1960, CLK => n4792, Q => 
                           RAM_1_121_port, QN => n_1163);
   RAM_reg_1_120_inst : DFFX1 port map( D => n1959, CLK => n4792, Q => 
                           RAM_1_120_port, QN => n_1164);
   RAM_reg_1_119_inst : DFFX1 port map( D => n1958, CLK => n4792, Q => 
                           RAM_1_119_port, QN => n_1165);
   RAM_reg_1_118_inst : DFFX1 port map( D => n1957, CLK => n4792, Q => 
                           RAM_1_118_port, QN => n_1166);
   RAM_reg_1_117_inst : DFFX1 port map( D => n1956, CLK => n4792, Q => 
                           RAM_1_117_port, QN => n_1167);
   RAM_reg_1_116_inst : DFFX1 port map( D => n1955, CLK => n4792, Q => 
                           RAM_1_116_port, QN => n_1168);
   RAM_reg_1_115_inst : DFFX1 port map( D => n1954, CLK => n4786, Q => 
                           RAM_1_115_port, QN => n_1169);
   RAM_reg_1_114_inst : DFFX1 port map( D => n1953, CLK => n4786, Q => 
                           RAM_1_114_port, QN => n_1170);
   RAM_reg_1_113_inst : DFFX1 port map( D => n1952, CLK => n4786, Q => 
                           RAM_1_113_port, QN => n_1171);
   RAM_reg_1_112_inst : DFFX1 port map( D => n1951, CLK => n4786, Q => 
                           RAM_1_112_port, QN => n_1172);
   RAM_reg_1_111_inst : DFFX1 port map( D => n1950, CLK => n4787, Q => 
                           RAM_1_111_port, QN => n_1173);
   RAM_reg_1_110_inst : DFFX1 port map( D => n1949, CLK => n4787, Q => 
                           RAM_1_110_port, QN => n_1174);
   RAM_reg_1_109_inst : DFFX1 port map( D => n1948, CLK => n4787, Q => 
                           RAM_1_109_port, QN => n_1175);
   RAM_reg_1_108_inst : DFFX1 port map( D => n1947, CLK => n4787, Q => 
                           RAM_1_108_port, QN => n_1176);
   RAM_reg_1_107_inst : DFFX1 port map( D => n1946, CLK => n4787, Q => 
                           RAM_1_107_port, QN => n_1177);
   RAM_reg_1_106_inst : DFFX1 port map( D => n1945, CLK => n4787, Q => 
                           RAM_1_106_port, QN => n_1178);
   RAM_reg_1_105_inst : DFFX1 port map( D => n1944, CLK => n4787, Q => 
                           RAM_1_105_port, QN => n_1179);
   RAM_reg_1_104_inst : DFFX1 port map( D => n1943, CLK => n4787, Q => 
                           RAM_1_104_port, QN => n_1180);
   RAM_reg_1_103_inst : DFFX1 port map( D => n1942, CLK => n4787, Q => 
                           RAM_1_103_port, QN => n_1181);
   RAM_reg_1_102_inst : DFFX1 port map( D => n1941, CLK => n4787, Q => 
                           RAM_1_102_port, QN => n_1182);
   RAM_reg_1_101_inst : DFFX1 port map( D => n1940, CLK => n4787, Q => 
                           RAM_1_101_port, QN => n_1183);
   RAM_reg_1_100_inst : DFFX1 port map( D => n1939, CLK => n4787, Q => 
                           RAM_1_100_port, QN => n_1184);
   RAM_reg_1_99_inst : DFFX1 port map( D => n1938, CLK => n4788, Q => 
                           RAM_1_99_port, QN => n_1185);
   RAM_reg_1_98_inst : DFFX1 port map( D => n1937, CLK => n4788, Q => 
                           RAM_1_98_port, QN => n_1186);
   RAM_reg_1_97_inst : DFFX1 port map( D => n1936, CLK => n4788, Q => 
                           RAM_1_97_port, QN => n_1187);
   RAM_reg_1_96_inst : DFFX1 port map( D => n1935, CLK => n4788, Q => 
                           RAM_1_96_port, QN => n_1188);
   RAM_reg_1_95_inst : DFFX1 port map( D => n1934, CLK => n4788, Q => 
                           RAM_1_95_port, QN => n_1189);
   RAM_reg_1_94_inst : DFFX1 port map( D => n1933, CLK => n4788, Q => 
                           RAM_1_94_port, QN => n_1190);
   RAM_reg_1_93_inst : DFFX1 port map( D => n1932, CLK => n4788, Q => 
                           RAM_1_93_port, QN => n_1191);
   RAM_reg_1_92_inst : DFFX1 port map( D => n1931, CLK => n4788, Q => 
                           RAM_1_92_port, QN => n_1192);
   RAM_reg_1_91_inst : DFFX1 port map( D => n1930, CLK => n4788, Q => 
                           RAM_1_91_port, QN => n_1193);
   RAM_reg_1_90_inst : DFFX1 port map( D => n1929, CLK => n4788, Q => 
                           RAM_1_90_port, QN => n_1194);
   RAM_reg_1_89_inst : DFFX1 port map( D => n1928, CLK => n4788, Q => 
                           RAM_1_89_port, QN => n_1195);
   RAM_reg_1_88_inst : DFFX1 port map( D => n1927, CLK => n4788, Q => 
                           RAM_1_88_port, QN => n_1196);
   RAM_reg_1_87_inst : DFFX1 port map( D => n1926, CLK => n4789, Q => 
                           RAM_1_87_port, QN => n_1197);
   RAM_reg_1_86_inst : DFFX1 port map( D => n1925, CLK => n4789, Q => 
                           RAM_1_86_port, QN => n_1198);
   RAM_reg_1_85_inst : DFFX1 port map( D => n1924, CLK => n4789, Q => 
                           RAM_1_85_port, QN => n_1199);
   RAM_reg_1_84_inst : DFFX1 port map( D => n1923, CLK => n4789, Q => 
                           RAM_1_84_port, QN => n_1200);
   RAM_reg_1_83_inst : DFFX1 port map( D => n1922, CLK => n4789, Q => 
                           RAM_1_83_port, QN => n_1201);
   RAM_reg_1_82_inst : DFFX1 port map( D => n1921, CLK => n4789, Q => 
                           RAM_1_82_port, QN => n_1202);
   RAM_reg_1_81_inst : DFFX1 port map( D => n1920, CLK => n4789, Q => 
                           RAM_1_81_port, QN => n_1203);
   RAM_reg_1_80_inst : DFFX1 port map( D => n1919, CLK => n4789, Q => 
                           RAM_1_80_port, QN => n_1204);
   RAM_reg_1_79_inst : DFFX1 port map( D => n1918, CLK => n4783, Q => 
                           RAM_1_79_port, QN => n_1205);
   RAM_reg_1_78_inst : DFFX1 port map( D => n1917, CLK => n4783, Q => 
                           RAM_1_78_port, QN => n_1206);
   RAM_reg_1_77_inst : DFFX1 port map( D => n1916, CLK => n4783, Q => 
                           RAM_1_77_port, QN => n_1207);
   RAM_reg_1_76_inst : DFFX1 port map( D => n1915, CLK => n4783, Q => 
                           RAM_1_76_port, QN => n_1208);
   RAM_reg_1_75_inst : DFFX1 port map( D => n1914, CLK => n4784, Q => 
                           RAM_1_75_port, QN => n_1209);
   RAM_reg_1_74_inst : DFFX1 port map( D => n1913, CLK => n4784, Q => 
                           RAM_1_74_port, QN => n_1210);
   RAM_reg_1_73_inst : DFFX1 port map( D => n1912, CLK => n4784, Q => 
                           RAM_1_73_port, QN => n_1211);
   RAM_reg_1_72_inst : DFFX1 port map( D => n1911, CLK => n4784, Q => 
                           RAM_1_72_port, QN => n_1212);
   RAM_reg_1_71_inst : DFFX1 port map( D => n1910, CLK => n4784, Q => 
                           RAM_1_71_port, QN => n_1213);
   RAM_reg_1_70_inst : DFFX1 port map( D => n1909, CLK => n4784, Q => 
                           RAM_1_70_port, QN => n_1214);
   RAM_reg_1_69_inst : DFFX1 port map( D => n1908, CLK => n4784, Q => 
                           RAM_1_69_port, QN => n_1215);
   RAM_reg_1_68_inst : DFFX1 port map( D => n1907, CLK => n4784, Q => 
                           RAM_1_68_port, QN => n_1216);
   RAM_reg_1_67_inst : DFFX1 port map( D => n1906, CLK => n4784, Q => 
                           RAM_1_67_port, QN => n_1217);
   RAM_reg_1_66_inst : DFFX1 port map( D => n1905, CLK => n4784, Q => 
                           RAM_1_66_port, QN => n_1218);
   RAM_reg_1_65_inst : DFFX1 port map( D => n1904, CLK => n4784, Q => 
                           RAM_1_65_port, QN => n_1219);
   RAM_reg_1_64_inst : DFFX1 port map( D => n1903, CLK => n4784, Q => 
                           RAM_1_64_port, QN => n_1220);
   RAM_reg_1_63_inst : DFFX1 port map( D => n1902, CLK => n4785, Q => 
                           RAM_1_63_port, QN => n_1221);
   RAM_reg_1_62_inst : DFFX1 port map( D => n1901, CLK => n4785, Q => 
                           RAM_1_62_port, QN => n_1222);
   RAM_reg_1_61_inst : DFFX1 port map( D => n1900, CLK => n4785, Q => 
                           RAM_1_61_port, QN => n_1223);
   RAM_reg_1_60_inst : DFFX1 port map( D => n1899, CLK => n4785, Q => 
                           RAM_1_60_port, QN => n_1224);
   RAM_reg_1_59_inst : DFFX1 port map( D => n1898, CLK => n4785, Q => 
                           RAM_1_59_port, QN => n_1225);
   RAM_reg_1_58_inst : DFFX1 port map( D => n1897, CLK => n4785, Q => 
                           RAM_1_58_port, QN => n_1226);
   RAM_reg_1_57_inst : DFFX1 port map( D => n1896, CLK => n4785, Q => 
                           RAM_1_57_port, QN => n_1227);
   RAM_reg_1_56_inst : DFFX1 port map( D => n1895, CLK => n4785, Q => 
                           RAM_1_56_port, QN => n_1228);
   RAM_reg_1_55_inst : DFFX1 port map( D => n1894, CLK => n4785, Q => 
                           RAM_1_55_port, QN => n_1229);
   RAM_reg_1_54_inst : DFFX1 port map( D => n1893, CLK => n4785, Q => 
                           RAM_1_54_port, QN => n_1230);
   RAM_reg_1_53_inst : DFFX1 port map( D => n1892, CLK => n4785, Q => 
                           RAM_1_53_port, QN => n_1231);
   RAM_reg_1_52_inst : DFFX1 port map( D => n1891, CLK => n4785, Q => 
                           RAM_1_52_port, QN => n_1232);
   RAM_reg_1_51_inst : DFFX1 port map( D => n1890, CLK => n4786, Q => 
                           RAM_1_51_port, QN => n_1233);
   RAM_reg_1_50_inst : DFFX1 port map( D => n1889, CLK => n4786, Q => 
                           RAM_1_50_port, QN => n_1234);
   RAM_reg_1_49_inst : DFFX1 port map( D => n1888, CLK => n4786, Q => 
                           RAM_1_49_port, QN => n_1235);
   RAM_reg_1_48_inst : DFFX1 port map( D => n1887, CLK => n4786, Q => 
                           RAM_1_48_port, QN => n_1236);
   RAM_reg_1_47_inst : DFFX1 port map( D => n1886, CLK => n4786, Q => 
                           RAM_1_47_port, QN => n_1237);
   RAM_reg_1_46_inst : DFFX1 port map( D => n1885, CLK => n4786, Q => 
                           RAM_1_46_port, QN => n_1238);
   RAM_reg_1_45_inst : DFFX1 port map( D => n1884, CLK => n4786, Q => 
                           RAM_1_45_port, QN => n_1239);
   RAM_reg_1_44_inst : DFFX1 port map( D => n1883, CLK => n4786, Q => 
                           RAM_1_44_port, QN => n_1240);
   RAM_reg_1_43_inst : DFFX1 port map( D => n1882, CLK => n4798, Q => 
                           RAM_1_43_port, QN => n_1241);
   RAM_reg_1_42_inst : DFFX1 port map( D => n1881, CLK => n4798, Q => 
                           RAM_1_42_port, QN => n_1242);
   RAM_reg_1_41_inst : DFFX1 port map( D => n1880, CLK => n4798, Q => 
                           RAM_1_41_port, QN => n_1243);
   RAM_reg_1_40_inst : DFFX1 port map( D => n1879, CLK => n4798, Q => 
                           RAM_1_40_port, QN => n_1244);
   RAM_reg_1_39_inst : DFFX1 port map( D => n1878, CLK => n4799, Q => 
                           RAM_1_39_port, QN => n_1245);
   RAM_reg_1_38_inst : DFFX1 port map( D => n1877, CLK => n4799, Q => 
                           RAM_1_38_port, QN => n_1246);
   RAM_reg_1_37_inst : DFFX1 port map( D => n1876, CLK => n4799, Q => 
                           RAM_1_37_port, QN => n_1247);
   RAM_reg_1_36_inst : DFFX1 port map( D => n1875, CLK => n4799, Q => 
                           RAM_1_36_port, QN => n_1248);
   RAM_reg_1_35_inst : DFFX1 port map( D => n1874, CLK => n4799, Q => 
                           RAM_1_35_port, QN => n_1249);
   RAM_reg_1_34_inst : DFFX1 port map( D => n1873, CLK => n4799, Q => 
                           RAM_1_34_port, QN => n_1250);
   RAM_reg_1_33_inst : DFFX1 port map( D => n1872, CLK => n4799, Q => 
                           RAM_1_33_port, QN => n_1251);
   RAM_reg_1_32_inst : DFFX1 port map( D => n1871, CLK => n4799, Q => 
                           RAM_1_32_port, QN => n_1252);
   RAM_reg_1_31_inst : DFFX1 port map( D => n1870, CLK => n4799, Q => 
                           RAM_1_31_port, QN => n_1253);
   RAM_reg_1_30_inst : DFFX1 port map( D => n1869, CLK => n4799, Q => 
                           RAM_1_30_port, QN => n_1254);
   RAM_reg_1_29_inst : DFFX1 port map( D => n1868, CLK => n4799, Q => 
                           RAM_1_29_port, QN => n_1255);
   RAM_reg_1_28_inst : DFFX1 port map( D => n1867, CLK => n4799, Q => 
                           RAM_1_28_port, QN => n_1256);
   RAM_reg_1_27_inst : DFFX1 port map( D => n1866, CLK => n4800, Q => 
                           RAM_1_27_port, QN => n_1257);
   RAM_reg_1_26_inst : DFFX1 port map( D => n1865, CLK => n4800, Q => 
                           RAM_1_26_port, QN => n_1258);
   RAM_reg_1_25_inst : DFFX1 port map( D => n1864, CLK => n4800, Q => 
                           RAM_1_25_port, QN => n_1259);
   RAM_reg_1_24_inst : DFFX1 port map( D => n1863, CLK => n4800, Q => 
                           RAM_1_24_port, QN => n_1260);
   RAM_reg_1_23_inst : DFFX1 port map( D => n1862, CLK => n4800, Q => 
                           RAM_1_23_port, QN => n_1261);
   RAM_reg_1_22_inst : DFFX1 port map( D => n1861, CLK => n4800, Q => 
                           RAM_1_22_port, QN => n_1262);
   RAM_reg_1_21_inst : DFFX1 port map( D => n1860, CLK => n4800, Q => 
                           RAM_1_21_port, QN => n_1263);
   RAM_reg_1_20_inst : DFFX1 port map( D => n1859, CLK => n4800, Q => 
                           RAM_1_20_port, QN => n_1264);
   RAM_reg_1_19_inst : DFFX1 port map( D => n1858, CLK => n4800, Q => 
                           RAM_1_19_port, QN => n_1265);
   RAM_reg_1_18_inst : DFFX1 port map( D => n1857, CLK => n4800, Q => 
                           RAM_1_18_port, QN => n_1266);
   RAM_reg_1_17_inst : DFFX1 port map( D => n1856, CLK => n4800, Q => 
                           RAM_1_17_port, QN => n_1267);
   RAM_reg_1_16_inst : DFFX1 port map( D => n1855, CLK => n4800, Q => 
                           RAM_1_16_port, QN => n_1268);
   RAM_reg_1_15_inst : DFFX1 port map( D => n1854, CLK => n4801, Q => 
                           RAM_1_15_port, QN => n_1269);
   RAM_reg_1_14_inst : DFFX1 port map( D => n1853, CLK => n4801, Q => 
                           RAM_1_14_port, QN => n_1270);
   RAM_reg_1_13_inst : DFFX1 port map( D => n1852, CLK => n4801, Q => 
                           RAM_1_13_port, QN => n_1271);
   RAM_reg_1_12_inst : DFFX1 port map( D => n1851, CLK => n4801, Q => 
                           RAM_1_12_port, QN => n_1272);
   RAM_reg_1_11_inst : DFFX1 port map( D => n1850, CLK => n4801, Q => 
                           RAM_1_11_port, QN => n_1273);
   RAM_reg_1_10_inst : DFFX1 port map( D => n1849, CLK => n4801, Q => 
                           RAM_1_10_port, QN => n_1274);
   RAM_reg_1_9_inst : DFFX1 port map( D => n1848, CLK => n4801, Q => 
                           RAM_1_9_port, QN => n_1275);
   RAM_reg_1_8_inst : DFFX1 port map( D => n1847, CLK => n4801, Q => 
                           RAM_1_8_port, QN => n_1276);
   RAM_reg_1_7_inst : DFFX1 port map( D => n1846, CLK => n4795, Q => 
                           RAM_1_7_port, QN => n_1277);
   RAM_reg_1_6_inst : DFFX1 port map( D => n1845, CLK => n4795, Q => 
                           RAM_1_6_port, QN => n_1278);
   RAM_reg_1_5_inst : DFFX1 port map( D => n1844, CLK => n4795, Q => 
                           RAM_1_5_port, QN => n_1279);
   RAM_reg_1_4_inst : DFFX1 port map( D => n1843, CLK => n4795, Q => 
                           RAM_1_4_port, QN => n_1280);
   RAM_reg_1_3_inst : DFFX1 port map( D => n1842, CLK => n4796, Q => 
                           RAM_1_3_port, QN => n_1281);
   RAM_reg_1_2_inst : DFFX1 port map( D => n1841, CLK => n4796, Q => 
                           RAM_1_2_port, QN => n_1282);
   RAM_reg_1_1_inst : DFFX1 port map( D => n1840, CLK => n4796, Q => 
                           RAM_1_1_port, QN => n_1283);
   RAM_reg_1_0_inst : DFFX1 port map( D => n1839, CLK => n4796, Q => 
                           RAM_1_0_port, QN => n_1284);
   RAM_reg_2_127_inst : DFFX1 port map( D => n1838, CLK => n4796, Q => 
                           RAM_2_127_port, QN => n_1285);
   RAM_reg_2_126_inst : DFFX1 port map( D => n1837, CLK => n4796, Q => 
                           RAM_2_126_port, QN => n_1286);
   RAM_reg_2_125_inst : DFFX1 port map( D => n1836, CLK => n4796, Q => 
                           RAM_2_125_port, QN => n_1287);
   RAM_reg_2_124_inst : DFFX1 port map( D => n1835, CLK => n4796, Q => 
                           RAM_2_124_port, QN => n_1288);
   RAM_reg_2_123_inst : DFFX1 port map( D => n1834, CLK => n4796, Q => 
                           RAM_2_123_port, QN => n_1289);
   RAM_reg_2_122_inst : DFFX1 port map( D => n1833, CLK => n4796, Q => 
                           RAM_2_122_port, QN => n_1290);
   RAM_reg_2_121_inst : DFFX1 port map( D => n1832, CLK => n4796, Q => 
                           RAM_2_121_port, QN => n_1291);
   RAM_reg_2_120_inst : DFFX1 port map( D => n1831, CLK => n4796, Q => 
                           RAM_2_120_port, QN => n_1292);
   RAM_reg_2_119_inst : DFFX1 port map( D => n1830, CLK => n4797, Q => 
                           RAM_2_119_port, QN => n_1293);
   RAM_reg_2_118_inst : DFFX1 port map( D => n1829, CLK => n4797, Q => 
                           RAM_2_118_port, QN => n_1294);
   RAM_reg_2_117_inst : DFFX1 port map( D => n1828, CLK => n4797, Q => 
                           RAM_2_117_port, QN => n_1295);
   RAM_reg_2_116_inst : DFFX1 port map( D => n1827, CLK => n4797, Q => 
                           RAM_2_116_port, QN => n_1296);
   RAM_reg_2_115_inst : DFFX1 port map( D => n1826, CLK => n4797, Q => 
                           RAM_2_115_port, QN => n_1297);
   RAM_reg_2_114_inst : DFFX1 port map( D => n1825, CLK => n4797, Q => 
                           RAM_2_114_port, QN => n_1298);
   RAM_reg_2_113_inst : DFFX1 port map( D => n1824, CLK => n4797, Q => 
                           RAM_2_113_port, QN => n_1299);
   RAM_reg_2_112_inst : DFFX1 port map( D => n1823, CLK => n4797, Q => 
                           RAM_2_112_port, QN => n_1300);
   RAM_reg_2_111_inst : DFFX1 port map( D => n1822, CLK => n4797, Q => 
                           RAM_2_111_port, QN => n_1301);
   RAM_reg_2_110_inst : DFFX1 port map( D => n1821, CLK => n4797, Q => 
                           RAM_2_110_port, QN => n_1302);
   RAM_reg_2_109_inst : DFFX1 port map( D => n1820, CLK => n4797, Q => 
                           RAM_2_109_port, QN => n_1303);
   RAM_reg_2_108_inst : DFFX1 port map( D => n1819, CLK => n4797, Q => 
                           RAM_2_108_port, QN => n_1304);
   RAM_reg_2_107_inst : DFFX1 port map( D => n1818, CLK => n4798, Q => 
                           RAM_2_107_port, QN => n_1305);
   RAM_reg_2_106_inst : DFFX1 port map( D => n1817, CLK => n4798, Q => 
                           RAM_2_106_port, QN => n_1306);
   RAM_reg_2_105_inst : DFFX1 port map( D => n1816, CLK => n4798, Q => 
                           RAM_2_105_port, QN => n_1307);
   RAM_reg_2_104_inst : DFFX1 port map( D => n1815, CLK => n4798, Q => 
                           RAM_2_104_port, QN => n_1308);
   RAM_reg_2_103_inst : DFFX1 port map( D => n1814, CLK => n4798, Q => 
                           RAM_2_103_port, QN => n_1309);
   RAM_reg_2_102_inst : DFFX1 port map( D => n1813, CLK => n4798, Q => 
                           RAM_2_102_port, QN => n_1310);
   RAM_reg_2_101_inst : DFFX1 port map( D => n1812, CLK => n4798, Q => 
                           RAM_2_101_port, QN => n_1311);
   RAM_reg_2_100_inst : DFFX1 port map( D => n1811, CLK => n4798, Q => 
                           RAM_2_100_port, QN => n_1312);
   RAM_reg_2_99_inst : DFFX1 port map( D => n1810, CLK => n4792, Q => 
                           RAM_2_99_port, QN => n_1313);
   RAM_reg_2_98_inst : DFFX1 port map( D => n1809, CLK => n4792, Q => 
                           RAM_2_98_port, QN => n_1314);
   RAM_reg_2_97_inst : DFFX1 port map( D => n1808, CLK => n4792, Q => 
                           RAM_2_97_port, QN => n_1315);
   RAM_reg_2_96_inst : DFFX1 port map( D => n1807, CLK => n4792, Q => 
                           RAM_2_96_port, QN => n_1316);
   RAM_reg_2_95_inst : DFFX1 port map( D => n1806, CLK => n4793, Q => 
                           RAM_2_95_port, QN => n_1317);
   RAM_reg_2_94_inst : DFFX1 port map( D => n1805, CLK => n4793, Q => 
                           RAM_2_94_port, QN => n_1318);
   RAM_reg_2_93_inst : DFFX1 port map( D => n1804, CLK => n4793, Q => 
                           RAM_2_93_port, QN => n_1319);
   RAM_reg_2_92_inst : DFFX1 port map( D => n1803, CLK => n4793, Q => 
                           RAM_2_92_port, QN => n_1320);
   RAM_reg_2_91_inst : DFFX1 port map( D => n1802, CLK => n4793, Q => 
                           RAM_2_91_port, QN => n_1321);
   RAM_reg_2_90_inst : DFFX1 port map( D => n1801, CLK => n4793, Q => 
                           RAM_2_90_port, QN => n_1322);
   RAM_reg_2_89_inst : DFFX1 port map( D => n1800, CLK => n4793, Q => 
                           RAM_2_89_port, QN => n_1323);
   RAM_reg_2_88_inst : DFFX1 port map( D => n1799, CLK => n4793, Q => 
                           RAM_2_88_port, QN => n_1324);
   RAM_reg_2_87_inst : DFFX1 port map( D => n1798, CLK => n4793, Q => 
                           RAM_2_87_port, QN => n_1325);
   RAM_reg_2_86_inst : DFFX1 port map( D => n1797, CLK => n4793, Q => 
                           RAM_2_86_port, QN => n_1326);
   RAM_reg_2_85_inst : DFFX1 port map( D => n1796, CLK => n4793, Q => 
                           RAM_2_85_port, QN => n_1327);
   RAM_reg_2_84_inst : DFFX1 port map( D => n1795, CLK => n4793, Q => 
                           RAM_2_84_port, QN => n_1328);
   RAM_reg_2_83_inst : DFFX1 port map( D => n1794, CLK => n4794, Q => 
                           RAM_2_83_port, QN => n_1329);
   RAM_reg_2_82_inst : DFFX1 port map( D => n1793, CLK => n4794, Q => 
                           RAM_2_82_port, QN => n_1330);
   RAM_reg_2_81_inst : DFFX1 port map( D => n1792, CLK => n4794, Q => 
                           RAM_2_81_port, QN => n_1331);
   RAM_reg_2_80_inst : DFFX1 port map( D => n1791, CLK => n4794, Q => 
                           RAM_2_80_port, QN => n_1332);
   RAM_reg_2_79_inst : DFFX1 port map( D => n1790, CLK => n4794, Q => 
                           RAM_2_79_port, QN => n_1333);
   RAM_reg_2_78_inst : DFFX1 port map( D => n1789, CLK => n4794, Q => 
                           RAM_2_78_port, QN => n_1334);
   RAM_reg_2_77_inst : DFFX1 port map( D => n1788, CLK => n4794, Q => 
                           RAM_2_77_port, QN => n_1335);
   RAM_reg_2_76_inst : DFFX1 port map( D => n1787, CLK => n4794, Q => 
                           RAM_2_76_port, QN => n_1336);
   RAM_reg_2_75_inst : DFFX1 port map( D => n1786, CLK => n4794, Q => 
                           RAM_2_75_port, QN => n_1337);
   RAM_reg_2_74_inst : DFFX1 port map( D => n1785, CLK => n4794, Q => 
                           RAM_2_74_port, QN => n_1338);
   RAM_reg_2_73_inst : DFFX1 port map( D => n1784, CLK => n4794, Q => 
                           RAM_2_73_port, QN => n_1339);
   RAM_reg_2_72_inst : DFFX1 port map( D => n1783, CLK => n4794, Q => 
                           RAM_2_72_port, QN => n_1340);
   RAM_reg_2_71_inst : DFFX1 port map( D => n1782, CLK => n4795, Q => 
                           RAM_2_71_port, QN => n_1341);
   RAM_reg_2_70_inst : DFFX1 port map( D => n1781, CLK => n4795, Q => 
                           RAM_2_70_port, QN => n_1342);
   RAM_reg_2_69_inst : DFFX1 port map( D => n1780, CLK => n4795, Q => 
                           RAM_2_69_port, QN => n_1343);
   RAM_reg_2_68_inst : DFFX1 port map( D => n1779, CLK => n4795, Q => 
                           RAM_2_68_port, QN => n_1344);
   RAM_reg_2_67_inst : DFFX1 port map( D => n1778, CLK => n4795, Q => 
                           RAM_2_67_port, QN => n_1345);
   RAM_reg_2_66_inst : DFFX1 port map( D => n1777, CLK => n4795, Q => 
                           RAM_2_66_port, QN => n_1346);
   RAM_reg_2_65_inst : DFFX1 port map( D => n1776, CLK => n4795, Q => 
                           RAM_2_65_port, QN => n_1347);
   RAM_reg_2_64_inst : DFFX1 port map( D => n1775, CLK => n4795, Q => 
                           RAM_2_64_port, QN => n_1348);
   RAM_reg_2_63_inst : DFFX1 port map( D => n1774, CLK => n4807, Q => 
                           RAM_2_63_port, QN => n_1349);
   RAM_reg_2_62_inst : DFFX1 port map( D => n1773, CLK => n4807, Q => 
                           RAM_2_62_port, QN => n_1350);
   RAM_reg_2_61_inst : DFFX1 port map( D => n1772, CLK => n4807, Q => 
                           RAM_2_61_port, QN => n_1351);
   RAM_reg_2_60_inst : DFFX1 port map( D => n1771, CLK => n4807, Q => 
                           RAM_2_60_port, QN => n_1352);
   RAM_reg_2_59_inst : DFFX1 port map( D => n1770, CLK => n4808, Q => 
                           RAM_2_59_port, QN => n_1353);
   RAM_reg_2_58_inst : DFFX1 port map( D => n1769, CLK => n4808, Q => 
                           RAM_2_58_port, QN => n_1354);
   RAM_reg_2_57_inst : DFFX1 port map( D => n1768, CLK => n4808, Q => 
                           RAM_2_57_port, QN => n_1355);
   RAM_reg_2_56_inst : DFFX1 port map( D => n1767, CLK => n4808, Q => 
                           RAM_2_56_port, QN => n_1356);
   RAM_reg_2_55_inst : DFFX1 port map( D => n1766, CLK => n4808, Q => 
                           RAM_2_55_port, QN => n_1357);
   RAM_reg_2_54_inst : DFFX1 port map( D => n1765, CLK => n4808, Q => 
                           RAM_2_54_port, QN => n_1358);
   RAM_reg_2_53_inst : DFFX1 port map( D => n1764, CLK => n4808, Q => 
                           RAM_2_53_port, QN => n_1359);
   RAM_reg_2_52_inst : DFFX1 port map( D => n1763, CLK => n4808, Q => 
                           RAM_2_52_port, QN => n_1360);
   RAM_reg_2_51_inst : DFFX1 port map( D => n1762, CLK => n4808, Q => 
                           RAM_2_51_port, QN => n_1361);
   RAM_reg_2_50_inst : DFFX1 port map( D => n1761, CLK => n4808, Q => 
                           RAM_2_50_port, QN => n_1362);
   RAM_reg_2_49_inst : DFFX1 port map( D => n1760, CLK => n4808, Q => 
                           RAM_2_49_port, QN => n_1363);
   RAM_reg_2_48_inst : DFFX1 port map( D => n1759, CLK => n4808, Q => 
                           RAM_2_48_port, QN => n_1364);
   RAM_reg_2_47_inst : DFFX1 port map( D => n1758, CLK => n4809, Q => 
                           RAM_2_47_port, QN => n_1365);
   RAM_reg_2_46_inst : DFFX1 port map( D => n1757, CLK => n4809, Q => 
                           RAM_2_46_port, QN => n_1366);
   RAM_reg_2_45_inst : DFFX1 port map( D => n1756, CLK => n4809, Q => 
                           RAM_2_45_port, QN => n_1367);
   RAM_reg_2_44_inst : DFFX1 port map( D => n1755, CLK => n4809, Q => 
                           RAM_2_44_port, QN => n_1368);
   RAM_reg_2_43_inst : DFFX1 port map( D => n1754, CLK => n4809, Q => 
                           RAM_2_43_port, QN => n_1369);
   RAM_reg_2_42_inst : DFFX1 port map( D => n1753, CLK => n4809, Q => 
                           RAM_2_42_port, QN => n_1370);
   RAM_reg_2_41_inst : DFFX1 port map( D => n1752, CLK => n4809, Q => 
                           RAM_2_41_port, QN => n_1371);
   RAM_reg_2_40_inst : DFFX1 port map( D => n1751, CLK => n4809, Q => 
                           RAM_2_40_port, QN => n_1372);
   RAM_reg_2_39_inst : DFFX1 port map( D => n1750, CLK => n4809, Q => 
                           RAM_2_39_port, QN => n_1373);
   RAM_reg_2_38_inst : DFFX1 port map( D => n1749, CLK => n4809, Q => 
                           RAM_2_38_port, QN => n_1374);
   RAM_reg_2_37_inst : DFFX1 port map( D => n1748, CLK => n4809, Q => 
                           RAM_2_37_port, QN => n_1375);
   RAM_reg_2_36_inst : DFFX1 port map( D => n1747, CLK => n4809, Q => 
                           RAM_2_36_port, QN => n_1376);
   RAM_reg_2_35_inst : DFFX1 port map( D => n1746, CLK => n4810, Q => 
                           RAM_2_35_port, QN => n_1377);
   RAM_reg_2_34_inst : DFFX1 port map( D => n1745, CLK => n4810, Q => 
                           RAM_2_34_port, QN => n_1378);
   RAM_reg_2_33_inst : DFFX1 port map( D => n1744, CLK => n4810, Q => 
                           RAM_2_33_port, QN => n_1379);
   RAM_reg_2_32_inst : DFFX1 port map( D => n1743, CLK => n4810, Q => 
                           RAM_2_32_port, QN => n_1380);
   RAM_reg_2_31_inst : DFFX1 port map( D => n1742, CLK => n4810, Q => 
                           RAM_2_31_port, QN => n_1381);
   RAM_reg_2_30_inst : DFFX1 port map( D => n1741, CLK => n4810, Q => 
                           RAM_2_30_port, QN => n_1382);
   RAM_reg_2_29_inst : DFFX1 port map( D => n1740, CLK => n4810, Q => 
                           RAM_2_29_port, QN => n_1383);
   RAM_reg_2_28_inst : DFFX1 port map( D => n1739, CLK => n4810, Q => 
                           RAM_2_28_port, QN => n_1384);
   RAM_reg_2_27_inst : DFFX1 port map( D => n1738, CLK => n4804, Q => 
                           RAM_2_27_port, QN => n_1385);
   RAM_reg_2_26_inst : DFFX1 port map( D => n1737, CLK => n4804, Q => 
                           RAM_2_26_port, QN => n_1386);
   RAM_reg_2_25_inst : DFFX1 port map( D => n1736, CLK => n4804, Q => 
                           RAM_2_25_port, QN => n_1387);
   RAM_reg_2_24_inst : DFFX1 port map( D => n1735, CLK => n4804, Q => 
                           RAM_2_24_port, QN => n_1388);
   RAM_reg_2_23_inst : DFFX1 port map( D => n1734, CLK => n4805, Q => 
                           RAM_2_23_port, QN => n_1389);
   RAM_reg_2_22_inst : DFFX1 port map( D => n1733, CLK => n4805, Q => 
                           RAM_2_22_port, QN => n_1390);
   RAM_reg_2_21_inst : DFFX1 port map( D => n1732, CLK => n4805, Q => 
                           RAM_2_21_port, QN => n_1391);
   RAM_reg_2_20_inst : DFFX1 port map( D => n1731, CLK => n4805, Q => 
                           RAM_2_20_port, QN => n_1392);
   RAM_reg_2_19_inst : DFFX1 port map( D => n1730, CLK => n4805, Q => 
                           RAM_2_19_port, QN => n_1393);
   RAM_reg_2_18_inst : DFFX1 port map( D => n1729, CLK => n4805, Q => 
                           RAM_2_18_port, QN => n_1394);
   RAM_reg_2_17_inst : DFFX1 port map( D => n1728, CLK => n4805, Q => 
                           RAM_2_17_port, QN => n_1395);
   RAM_reg_2_16_inst : DFFX1 port map( D => n1727, CLK => n4805, Q => 
                           RAM_2_16_port, QN => n_1396);
   RAM_reg_2_15_inst : DFFX1 port map( D => n1726, CLK => n4805, Q => 
                           RAM_2_15_port, QN => n_1397);
   RAM_reg_2_14_inst : DFFX1 port map( D => n1725, CLK => n4805, Q => 
                           RAM_2_14_port, QN => n_1398);
   RAM_reg_2_13_inst : DFFX1 port map( D => n1724, CLK => n4805, Q => 
                           RAM_2_13_port, QN => n_1399);
   RAM_reg_2_12_inst : DFFX1 port map( D => n1723, CLK => n4805, Q => 
                           RAM_2_12_port, QN => n_1400);
   RAM_reg_2_11_inst : DFFX1 port map( D => n1722, CLK => n4806, Q => 
                           RAM_2_11_port, QN => n_1401);
   RAM_reg_2_10_inst : DFFX1 port map( D => n1721, CLK => n4806, Q => 
                           RAM_2_10_port, QN => n_1402);
   RAM_reg_2_9_inst : DFFX1 port map( D => n1720, CLK => n4806, Q => 
                           RAM_2_9_port, QN => n_1403);
   RAM_reg_2_8_inst : DFFX1 port map( D => n1719, CLK => n4806, Q => 
                           RAM_2_8_port, QN => n_1404);
   RAM_reg_2_7_inst : DFFX1 port map( D => n1718, CLK => n4806, Q => 
                           RAM_2_7_port, QN => n_1405);
   RAM_reg_2_6_inst : DFFX1 port map( D => n1717, CLK => n4806, Q => 
                           RAM_2_6_port, QN => n_1406);
   RAM_reg_2_5_inst : DFFX1 port map( D => n1716, CLK => n4806, Q => 
                           RAM_2_5_port, QN => n_1407);
   RAM_reg_2_4_inst : DFFX1 port map( D => n1715, CLK => n4806, Q => 
                           RAM_2_4_port, QN => n_1408);
   RAM_reg_2_3_inst : DFFX1 port map( D => n1714, CLK => n4806, Q => 
                           RAM_2_3_port, QN => n_1409);
   RAM_reg_2_2_inst : DFFX1 port map( D => n1713, CLK => n4806, Q => 
                           RAM_2_2_port, QN => n_1410);
   RAM_reg_2_1_inst : DFFX1 port map( D => n1712, CLK => n4806, Q => 
                           RAM_2_1_port, QN => n_1411);
   RAM_reg_2_0_inst : DFFX1 port map( D => n1711, CLK => n4806, Q => 
                           RAM_2_0_port, QN => n_1412);
   RAM_reg_3_127_inst : DFFX1 port map( D => n1710, CLK => n4807, Q => 
                           RAM_3_127_port, QN => n_1413);
   RAM_reg_3_126_inst : DFFX1 port map( D => n1709, CLK => n4807, Q => 
                           RAM_3_126_port, QN => n_1414);
   RAM_reg_3_125_inst : DFFX1 port map( D => n1708, CLK => n4807, Q => 
                           RAM_3_125_port, QN => n_1415);
   RAM_reg_3_124_inst : DFFX1 port map( D => n1707, CLK => n4807, Q => 
                           RAM_3_124_port, QN => n_1416);
   RAM_reg_3_123_inst : DFFX1 port map( D => n1706, CLK => n4807, Q => 
                           RAM_3_123_port, QN => n_1417);
   RAM_reg_3_122_inst : DFFX1 port map( D => n1705, CLK => n4807, Q => 
                           RAM_3_122_port, QN => n_1418);
   RAM_reg_3_121_inst : DFFX1 port map( D => n1704, CLK => n4807, Q => 
                           RAM_3_121_port, QN => n_1419);
   RAM_reg_3_120_inst : DFFX1 port map( D => n1703, CLK => n4807, Q => 
                           RAM_3_120_port, QN => n_1420);
   RAM_reg_3_119_inst : DFFX1 port map( D => n1702, CLK => n4801, Q => 
                           RAM_3_119_port, QN => n_1421);
   RAM_reg_3_118_inst : DFFX1 port map( D => n1701, CLK => n4801, Q => 
                           RAM_3_118_port, QN => n_1422);
   RAM_reg_3_117_inst : DFFX1 port map( D => n1700, CLK => n4801, Q => 
                           RAM_3_117_port, QN => n_1423);
   RAM_reg_3_116_inst : DFFX1 port map( D => n1699, CLK => n4801, Q => 
                           RAM_3_116_port, QN => n_1424);
   RAM_reg_3_115_inst : DFFX1 port map( D => n1698, CLK => n4802, Q => 
                           RAM_3_115_port, QN => n_1425);
   RAM_reg_3_114_inst : DFFX1 port map( D => n1697, CLK => n4802, Q => 
                           RAM_3_114_port, QN => n_1426);
   RAM_reg_3_113_inst : DFFX1 port map( D => n1696, CLK => n4802, Q => 
                           RAM_3_113_port, QN => n_1427);
   RAM_reg_3_112_inst : DFFX1 port map( D => n1695, CLK => n4802, Q => 
                           RAM_3_112_port, QN => n_1428);
   RAM_reg_3_111_inst : DFFX1 port map( D => n1694, CLK => n4802, Q => 
                           RAM_3_111_port, QN => n_1429);
   RAM_reg_3_110_inst : DFFX1 port map( D => n1693, CLK => n4802, Q => 
                           RAM_3_110_port, QN => n_1430);
   RAM_reg_3_109_inst : DFFX1 port map( D => n1692, CLK => n4802, Q => 
                           RAM_3_109_port, QN => n_1431);
   RAM_reg_3_108_inst : DFFX1 port map( D => n1691, CLK => n4802, Q => 
                           RAM_3_108_port, QN => n_1432);
   RAM_reg_3_107_inst : DFFX1 port map( D => n1690, CLK => n4802, Q => 
                           RAM_3_107_port, QN => n_1433);
   RAM_reg_3_106_inst : DFFX1 port map( D => n1689, CLK => n4802, Q => 
                           RAM_3_106_port, QN => n_1434);
   RAM_reg_3_105_inst : DFFX1 port map( D => n1688, CLK => n4802, Q => 
                           RAM_3_105_port, QN => n_1435);
   RAM_reg_3_104_inst : DFFX1 port map( D => n1687, CLK => n4802, Q => 
                           RAM_3_104_port, QN => n_1436);
   RAM_reg_3_103_inst : DFFX1 port map( D => n1686, CLK => n4803, Q => 
                           RAM_3_103_port, QN => n_1437);
   RAM_reg_3_102_inst : DFFX1 port map( D => n1685, CLK => n4803, Q => 
                           RAM_3_102_port, QN => n_1438);
   RAM_reg_3_101_inst : DFFX1 port map( D => n1684, CLK => n4803, Q => 
                           RAM_3_101_port, QN => n_1439);
   RAM_reg_3_100_inst : DFFX1 port map( D => n1683, CLK => n4803, Q => 
                           RAM_3_100_port, QN => n_1440);
   RAM_reg_3_99_inst : DFFX1 port map( D => n1682, CLK => n4803, Q => 
                           RAM_3_99_port, QN => n_1441);
   RAM_reg_3_98_inst : DFFX1 port map( D => n1681, CLK => n4803, Q => 
                           RAM_3_98_port, QN => n_1442);
   RAM_reg_3_97_inst : DFFX1 port map( D => n1680, CLK => n4803, Q => 
                           RAM_3_97_port, QN => n_1443);
   RAM_reg_3_96_inst : DFFX1 port map( D => n1679, CLK => n4803, Q => 
                           RAM_3_96_port, QN => n_1444);
   RAM_reg_3_95_inst : DFFX1 port map( D => n1678, CLK => n4803, Q => 
                           RAM_3_95_port, QN => n_1445);
   RAM_reg_3_94_inst : DFFX1 port map( D => n1677, CLK => n4803, Q => 
                           RAM_3_94_port, QN => n_1446);
   RAM_reg_3_93_inst : DFFX1 port map( D => n1676, CLK => n4803, Q => 
                           RAM_3_93_port, QN => n_1447);
   RAM_reg_3_92_inst : DFFX1 port map( D => n1675, CLK => n4803, Q => 
                           RAM_3_92_port, QN => n_1448);
   RAM_reg_3_91_inst : DFFX1 port map( D => n1674, CLK => n4804, Q => 
                           RAM_3_91_port, QN => n_1449);
   RAM_reg_3_90_inst : DFFX1 port map( D => n1673, CLK => n4804, Q => 
                           RAM_3_90_port, QN => n_1450);
   RAM_reg_3_89_inst : DFFX1 port map( D => n1672, CLK => n4804, Q => 
                           RAM_3_89_port, QN => n_1451);
   RAM_reg_3_88_inst : DFFX1 port map( D => n1671, CLK => n4804, Q => 
                           RAM_3_88_port, QN => n_1452);
   RAM_reg_3_87_inst : DFFX1 port map( D => n1670, CLK => n4804, Q => 
                           RAM_3_87_port, QN => n_1453);
   RAM_reg_3_86_inst : DFFX1 port map( D => n1669, CLK => n4804, Q => 
                           RAM_3_86_port, QN => n_1454);
   RAM_reg_3_85_inst : DFFX1 port map( D => n1668, CLK => n4804, Q => 
                           RAM_3_85_port, QN => n_1455);
   RAM_reg_3_84_inst : DFFX1 port map( D => n1667, CLK => n4804, Q => 
                           RAM_3_84_port, QN => n_1456);
   RAM_reg_3_83_inst : DFFX1 port map( D => n1666, CLK => n4816, Q => 
                           RAM_3_83_port, QN => n_1457);
   RAM_reg_3_82_inst : DFFX1 port map( D => n1665, CLK => n4816, Q => 
                           RAM_3_82_port, QN => n_1458);
   RAM_reg_3_81_inst : DFFX1 port map( D => n1664, CLK => n4816, Q => 
                           RAM_3_81_port, QN => n_1459);
   RAM_reg_3_80_inst : DFFX1 port map( D => n1663, CLK => n4816, Q => 
                           RAM_3_80_port, QN => n_1460);
   RAM_reg_3_79_inst : DFFX1 port map( D => n1662, CLK => n4817, Q => 
                           RAM_3_79_port, QN => n_1461);
   RAM_reg_3_78_inst : DFFX1 port map( D => n1661, CLK => n4817, Q => 
                           RAM_3_78_port, QN => n_1462);
   RAM_reg_3_77_inst : DFFX1 port map( D => n1660, CLK => n4817, Q => 
                           RAM_3_77_port, QN => n_1463);
   RAM_reg_3_76_inst : DFFX1 port map( D => n1659, CLK => n4817, Q => 
                           RAM_3_76_port, QN => n_1464);
   RAM_reg_3_75_inst : DFFX1 port map( D => n1658, CLK => n4817, Q => 
                           RAM_3_75_port, QN => n_1465);
   RAM_reg_3_74_inst : DFFX1 port map( D => n1657, CLK => n4817, Q => 
                           RAM_3_74_port, QN => n_1466);
   RAM_reg_3_73_inst : DFFX1 port map( D => n1656, CLK => n4817, Q => 
                           RAM_3_73_port, QN => n_1467);
   RAM_reg_3_72_inst : DFFX1 port map( D => n1655, CLK => n4817, Q => 
                           RAM_3_72_port, QN => n_1468);
   RAM_reg_3_71_inst : DFFX1 port map( D => n1654, CLK => n4817, Q => 
                           RAM_3_71_port, QN => n_1469);
   RAM_reg_3_70_inst : DFFX1 port map( D => n1653, CLK => n4817, Q => 
                           RAM_3_70_port, QN => n_1470);
   RAM_reg_3_69_inst : DFFX1 port map( D => n1652, CLK => n4817, Q => 
                           RAM_3_69_port, QN => n_1471);
   RAM_reg_3_68_inst : DFFX1 port map( D => n1651, CLK => n4817, Q => 
                           RAM_3_68_port, QN => n_1472);
   RAM_reg_3_67_inst : DFFX1 port map( D => n1650, CLK => n4818, Q => 
                           RAM_3_67_port, QN => n_1473);
   RAM_reg_3_66_inst : DFFX1 port map( D => n1649, CLK => n4818, Q => 
                           RAM_3_66_port, QN => n_1474);
   RAM_reg_3_65_inst : DFFX1 port map( D => n1648, CLK => n4818, Q => 
                           RAM_3_65_port, QN => n_1475);
   RAM_reg_3_64_inst : DFFX1 port map( D => n1647, CLK => n4818, Q => 
                           RAM_3_64_port, QN => n_1476);
   RAM_reg_3_63_inst : DFFX1 port map( D => n1646, CLK => n4818, Q => 
                           RAM_3_63_port, QN => n_1477);
   RAM_reg_3_62_inst : DFFX1 port map( D => n1645, CLK => n4818, Q => 
                           RAM_3_62_port, QN => n_1478);
   RAM_reg_3_61_inst : DFFX1 port map( D => n1644, CLK => n4818, Q => 
                           RAM_3_61_port, QN => n_1479);
   RAM_reg_3_60_inst : DFFX1 port map( D => n1643, CLK => n4818, Q => 
                           RAM_3_60_port, QN => n_1480);
   RAM_reg_3_59_inst : DFFX1 port map( D => n1642, CLK => n4818, Q => 
                           RAM_3_59_port, QN => n_1481);
   RAM_reg_3_58_inst : DFFX1 port map( D => n1641, CLK => n4818, Q => 
                           RAM_3_58_port, QN => n_1482);
   RAM_reg_3_57_inst : DFFX1 port map( D => n1640, CLK => n4818, Q => 
                           RAM_3_57_port, QN => n_1483);
   RAM_reg_3_56_inst : DFFX1 port map( D => n1639, CLK => n4818, Q => 
                           RAM_3_56_port, QN => n_1484);
   RAM_reg_3_55_inst : DFFX1 port map( D => n1638, CLK => n4819, Q => 
                           RAM_3_55_port, QN => n_1485);
   RAM_reg_3_54_inst : DFFX1 port map( D => n1637, CLK => n4819, Q => 
                           RAM_3_54_port, QN => n_1486);
   RAM_reg_3_53_inst : DFFX1 port map( D => n1636, CLK => n4819, Q => 
                           RAM_3_53_port, QN => n_1487);
   RAM_reg_3_52_inst : DFFX1 port map( D => n1635, CLK => n4819, Q => 
                           RAM_3_52_port, QN => n_1488);
   RAM_reg_3_51_inst : DFFX1 port map( D => n1634, CLK => n4819, Q => 
                           RAM_3_51_port, QN => n_1489);
   RAM_reg_3_50_inst : DFFX1 port map( D => n1633, CLK => n4819, Q => 
                           RAM_3_50_port, QN => n_1490);
   RAM_reg_3_49_inst : DFFX1 port map( D => n1632, CLK => n4819, Q => 
                           RAM_3_49_port, QN => n_1491);
   RAM_reg_3_48_inst : DFFX1 port map( D => n1631, CLK => n4819, Q => 
                           RAM_3_48_port, QN => n_1492);
   RAM_reg_3_47_inst : DFFX1 port map( D => n1630, CLK => n4813, Q => 
                           RAM_3_47_port, QN => n_1493);
   RAM_reg_3_46_inst : DFFX1 port map( D => n1629, CLK => n4813, Q => 
                           RAM_3_46_port, QN => n_1494);
   RAM_reg_3_45_inst : DFFX1 port map( D => n1628, CLK => n4813, Q => 
                           RAM_3_45_port, QN => n_1495);
   RAM_reg_3_44_inst : DFFX1 port map( D => n1627, CLK => n4813, Q => 
                           RAM_3_44_port, QN => n_1496);
   RAM_reg_3_43_inst : DFFX1 port map( D => n1626, CLK => n4814, Q => 
                           RAM_3_43_port, QN => n_1497);
   RAM_reg_3_42_inst : DFFX1 port map( D => n1625, CLK => n4814, Q => 
                           RAM_3_42_port, QN => n_1498);
   RAM_reg_3_41_inst : DFFX1 port map( D => n1624, CLK => n4814, Q => 
                           RAM_3_41_port, QN => n_1499);
   RAM_reg_3_40_inst : DFFX1 port map( D => n1623, CLK => n4814, Q => 
                           RAM_3_40_port, QN => n_1500);
   RAM_reg_3_39_inst : DFFX1 port map( D => n1622, CLK => n4814, Q => 
                           RAM_3_39_port, QN => n_1501);
   RAM_reg_3_38_inst : DFFX1 port map( D => n1621, CLK => n4814, Q => 
                           RAM_3_38_port, QN => n_1502);
   RAM_reg_3_37_inst : DFFX1 port map( D => n1620, CLK => n4814, Q => 
                           RAM_3_37_port, QN => n_1503);
   RAM_reg_3_36_inst : DFFX1 port map( D => n1619, CLK => n4814, Q => 
                           RAM_3_36_port, QN => n_1504);
   RAM_reg_3_35_inst : DFFX1 port map( D => n1618, CLK => n4814, Q => 
                           RAM_3_35_port, QN => n_1505);
   RAM_reg_3_34_inst : DFFX1 port map( D => n1617, CLK => n4814, Q => 
                           RAM_3_34_port, QN => n_1506);
   RAM_reg_3_33_inst : DFFX1 port map( D => n1616, CLK => n4814, Q => 
                           RAM_3_33_port, QN => n_1507);
   RAM_reg_3_32_inst : DFFX1 port map( D => n1615, CLK => n4814, Q => 
                           RAM_3_32_port, QN => n_1508);
   RAM_reg_3_31_inst : DFFX1 port map( D => n1614, CLK => n4815, Q => 
                           RAM_3_31_port, QN => n_1509);
   RAM_reg_3_30_inst : DFFX1 port map( D => n1613, CLK => n4815, Q => 
                           RAM_3_30_port, QN => n_1510);
   RAM_reg_3_29_inst : DFFX1 port map( D => n1612, CLK => n4815, Q => 
                           RAM_3_29_port, QN => n_1511);
   RAM_reg_3_28_inst : DFFX1 port map( D => n1611, CLK => n4815, Q => 
                           RAM_3_28_port, QN => n_1512);
   RAM_reg_3_27_inst : DFFX1 port map( D => n1610, CLK => n4815, Q => 
                           RAM_3_27_port, QN => n_1513);
   RAM_reg_3_26_inst : DFFX1 port map( D => n1609, CLK => n4815, Q => 
                           RAM_3_26_port, QN => n_1514);
   RAM_reg_3_25_inst : DFFX1 port map( D => n1608, CLK => n4815, Q => 
                           RAM_3_25_port, QN => n_1515);
   RAM_reg_3_24_inst : DFFX1 port map( D => n1607, CLK => n4815, Q => 
                           RAM_3_24_port, QN => n_1516);
   RAM_reg_3_23_inst : DFFX1 port map( D => n1606, CLK => n4815, Q => 
                           RAM_3_23_port, QN => n_1517);
   RAM_reg_3_22_inst : DFFX1 port map( D => n1605, CLK => n4815, Q => 
                           RAM_3_22_port, QN => n_1518);
   RAM_reg_3_21_inst : DFFX1 port map( D => n1604, CLK => n4815, Q => 
                           RAM_3_21_port, QN => n_1519);
   RAM_reg_3_20_inst : DFFX1 port map( D => n1603, CLK => n4815, Q => 
                           RAM_3_20_port, QN => n_1520);
   RAM_reg_3_19_inst : DFFX1 port map( D => n1602, CLK => n4816, Q => 
                           RAM_3_19_port, QN => n_1521);
   RAM_reg_3_18_inst : DFFX1 port map( D => n1601, CLK => n4816, Q => 
                           RAM_3_18_port, QN => n_1522);
   RAM_reg_3_17_inst : DFFX1 port map( D => n1600, CLK => n4816, Q => 
                           RAM_3_17_port, QN => n_1523);
   RAM_reg_3_16_inst : DFFX1 port map( D => n1599, CLK => n4816, Q => 
                           RAM_3_16_port, QN => n_1524);
   RAM_reg_3_15_inst : DFFX1 port map( D => n1598, CLK => n4816, Q => 
                           RAM_3_15_port, QN => n_1525);
   RAM_reg_3_14_inst : DFFX1 port map( D => n1597, CLK => n4816, Q => 
                           RAM_3_14_port, QN => n_1526);
   RAM_reg_3_13_inst : DFFX1 port map( D => n1596, CLK => n4816, Q => 
                           RAM_3_13_port, QN => n_1527);
   RAM_reg_3_12_inst : DFFX1 port map( D => n1595, CLK => n4816, Q => 
                           RAM_3_12_port, QN => n_1528);
   RAM_reg_3_11_inst : DFFX1 port map( D => n1594, CLK => n4810, Q => 
                           RAM_3_11_port, QN => n_1529);
   RAM_reg_3_10_inst : DFFX1 port map( D => n1593, CLK => n4810, Q => 
                           RAM_3_10_port, QN => n_1530);
   RAM_reg_3_9_inst : DFFX1 port map( D => n1592, CLK => n4810, Q => 
                           RAM_3_9_port, QN => n_1531);
   RAM_reg_3_8_inst : DFFX1 port map( D => n1591, CLK => n4810, Q => 
                           RAM_3_8_port, QN => n_1532);
   RAM_reg_3_7_inst : DFFX1 port map( D => n1590, CLK => n4811, Q => 
                           RAM_3_7_port, QN => n_1533);
   RAM_reg_3_6_inst : DFFX1 port map( D => n1589, CLK => n4811, Q => 
                           RAM_3_6_port, QN => n_1534);
   RAM_reg_3_5_inst : DFFX1 port map( D => n1588, CLK => n4811, Q => 
                           RAM_3_5_port, QN => n_1535);
   RAM_reg_3_4_inst : DFFX1 port map( D => n1587, CLK => n4811, Q => 
                           RAM_3_4_port, QN => n_1536);
   RAM_reg_3_3_inst : DFFX1 port map( D => n1586, CLK => n4811, Q => 
                           RAM_3_3_port, QN => n_1537);
   RAM_reg_3_2_inst : DFFX1 port map( D => n1585, CLK => n4811, Q => 
                           RAM_3_2_port, QN => n_1538);
   RAM_reg_3_1_inst : DFFX1 port map( D => n1584, CLK => n4811, Q => 
                           RAM_3_1_port, QN => n_1539);
   RAM_reg_3_0_inst : DFFX1 port map( D => n1583, CLK => n4811, Q => 
                           RAM_3_0_port, QN => n_1540);
   RAM_reg_4_127_inst : DFFX1 port map( D => n1582, CLK => n4811, Q => 
                           RAM_4_127_port, QN => n_1541);
   RAM_reg_4_126_inst : DFFX1 port map( D => n1581, CLK => n4811, Q => 
                           RAM_4_126_port, QN => n_1542);
   RAM_reg_4_125_inst : DFFX1 port map( D => n1580, CLK => n4811, Q => 
                           RAM_4_125_port, QN => n_1543);
   RAM_reg_4_124_inst : DFFX1 port map( D => n1579, CLK => n4811, Q => 
                           RAM_4_124_port, QN => n_1544);
   RAM_reg_4_123_inst : DFFX1 port map( D => n1578, CLK => n4812, Q => 
                           RAM_4_123_port, QN => n_1545);
   RAM_reg_4_122_inst : DFFX1 port map( D => n1577, CLK => n4812, Q => 
                           RAM_4_122_port, QN => n_1546);
   RAM_reg_4_121_inst : DFFX1 port map( D => n1576, CLK => n4812, Q => 
                           RAM_4_121_port, QN => n_1547);
   RAM_reg_4_120_inst : DFFX1 port map( D => n1575, CLK => n4812, Q => 
                           RAM_4_120_port, QN => n_1548);
   RAM_reg_4_119_inst : DFFX1 port map( D => n1574, CLK => n4812, Q => 
                           RAM_4_119_port, QN => n_1549);
   RAM_reg_4_118_inst : DFFX1 port map( D => n1573, CLK => n4812, Q => 
                           RAM_4_118_port, QN => n_1550);
   RAM_reg_4_117_inst : DFFX1 port map( D => n1572, CLK => n4812, Q => 
                           RAM_4_117_port, QN => n_1551);
   RAM_reg_4_116_inst : DFFX1 port map( D => n1571, CLK => n4812, Q => 
                           RAM_4_116_port, QN => n_1552);
   RAM_reg_4_115_inst : DFFX1 port map( D => n1570, CLK => n4812, Q => 
                           RAM_4_115_port, QN => n_1553);
   RAM_reg_4_114_inst : DFFX1 port map( D => n1569, CLK => n4812, Q => 
                           RAM_4_114_port, QN => n_1554);
   RAM_reg_4_113_inst : DFFX1 port map( D => n1568, CLK => n4812, Q => 
                           RAM_4_113_port, QN => n_1555);
   RAM_reg_4_112_inst : DFFX1 port map( D => n1567, CLK => n4812, Q => 
                           RAM_4_112_port, QN => n_1556);
   RAM_reg_4_111_inst : DFFX1 port map( D => n1566, CLK => n4813, Q => 
                           RAM_4_111_port, QN => n_1557);
   RAM_reg_4_110_inst : DFFX1 port map( D => n1565, CLK => n4813, Q => 
                           RAM_4_110_port, QN => n_1558);
   RAM_reg_4_109_inst : DFFX1 port map( D => n1564, CLK => n4813, Q => 
                           RAM_4_109_port, QN => n_1559);
   RAM_reg_4_108_inst : DFFX1 port map( D => n1563, CLK => n4813, Q => 
                           RAM_4_108_port, QN => n_1560);
   RAM_reg_4_107_inst : DFFX1 port map( D => n1562, CLK => n4813, Q => 
                           RAM_4_107_port, QN => n_1561);
   RAM_reg_4_106_inst : DFFX1 port map( D => n1561, CLK => n4813, Q => 
                           RAM_4_106_port, QN => n_1562);
   RAM_reg_4_105_inst : DFFX1 port map( D => n1560, CLK => n4813, Q => 
                           RAM_4_105_port, QN => n_1563);
   RAM_reg_4_104_inst : DFFX1 port map( D => n1559, CLK => n4813, Q => 
                           RAM_4_104_port, QN => n_1564);
   RAM_reg_4_103_inst : DFFX1 port map( D => n1558, CLK => n4825, Q => 
                           RAM_4_103_port, QN => n_1565);
   RAM_reg_4_102_inst : DFFX1 port map( D => n1557, CLK => n4825, Q => 
                           RAM_4_102_port, QN => n_1566);
   RAM_reg_4_101_inst : DFFX1 port map( D => n1556, CLK => n4825, Q => 
                           RAM_4_101_port, QN => n_1567);
   RAM_reg_4_100_inst : DFFX1 port map( D => n1555, CLK => n4825, Q => 
                           RAM_4_100_port, QN => n_1568);
   RAM_reg_4_99_inst : DFFX1 port map( D => n1554, CLK => n4826, Q => 
                           RAM_4_99_port, QN => n_1569);
   RAM_reg_4_98_inst : DFFX1 port map( D => n1553, CLK => n4826, Q => 
                           RAM_4_98_port, QN => n_1570);
   RAM_reg_4_97_inst : DFFX1 port map( D => n1552, CLK => n4826, Q => 
                           RAM_4_97_port, QN => n_1571);
   RAM_reg_4_96_inst : DFFX1 port map( D => n1551, CLK => n4826, Q => 
                           RAM_4_96_port, QN => n_1572);
   RAM_reg_4_95_inst : DFFX1 port map( D => n1550, CLK => n4826, Q => 
                           RAM_4_95_port, QN => n_1573);
   RAM_reg_4_94_inst : DFFX1 port map( D => n1549, CLK => n4826, Q => 
                           RAM_4_94_port, QN => n_1574);
   RAM_reg_4_93_inst : DFFX1 port map( D => n1548, CLK => n4826, Q => 
                           RAM_4_93_port, QN => n_1575);
   RAM_reg_4_92_inst : DFFX1 port map( D => n1547, CLK => n4826, Q => 
                           RAM_4_92_port, QN => n_1576);
   RAM_reg_4_91_inst : DFFX1 port map( D => n1546, CLK => n4826, Q => 
                           RAM_4_91_port, QN => n_1577);
   RAM_reg_4_90_inst : DFFX1 port map( D => n1545, CLK => n4826, Q => 
                           RAM_4_90_port, QN => n_1578);
   RAM_reg_4_89_inst : DFFX1 port map( D => n1544, CLK => n4826, Q => 
                           RAM_4_89_port, QN => n_1579);
   RAM_reg_4_88_inst : DFFX1 port map( D => n1543, CLK => n4826, Q => 
                           RAM_4_88_port, QN => n_1580);
   RAM_reg_4_87_inst : DFFX1 port map( D => n1542, CLK => n4827, Q => 
                           RAM_4_87_port, QN => n_1581);
   RAM_reg_4_86_inst : DFFX1 port map( D => n1541, CLK => n4827, Q => 
                           RAM_4_86_port, QN => n_1582);
   RAM_reg_4_85_inst : DFFX1 port map( D => n1540, CLK => n4827, Q => 
                           RAM_4_85_port, QN => n_1583);
   RAM_reg_4_84_inst : DFFX1 port map( D => n1539, CLK => n4827, Q => 
                           RAM_4_84_port, QN => n_1584);
   RAM_reg_4_83_inst : DFFX1 port map( D => n1538, CLK => n4827, Q => 
                           RAM_4_83_port, QN => n_1585);
   RAM_reg_4_82_inst : DFFX1 port map( D => n1537, CLK => n4827, Q => 
                           RAM_4_82_port, QN => n_1586);
   RAM_reg_4_81_inst : DFFX1 port map( D => n1536, CLK => n4827, Q => 
                           RAM_4_81_port, QN => n_1587);
   RAM_reg_4_80_inst : DFFX1 port map( D => n1535, CLK => n4827, Q => 
                           RAM_4_80_port, QN => n_1588);
   RAM_reg_4_79_inst : DFFX1 port map( D => n1534, CLK => n4827, Q => 
                           RAM_4_79_port, QN => n_1589);
   RAM_reg_4_78_inst : DFFX1 port map( D => n1533, CLK => n4827, Q => 
                           RAM_4_78_port, QN => n_1590);
   RAM_reg_4_77_inst : DFFX1 port map( D => n1532, CLK => n4827, Q => 
                           RAM_4_77_port, QN => n_1591);
   RAM_reg_4_76_inst : DFFX1 port map( D => n1531, CLK => n4827, Q => 
                           RAM_4_76_port, QN => n_1592);
   RAM_reg_4_75_inst : DFFX1 port map( D => n1530, CLK => n4828, Q => 
                           RAM_4_75_port, QN => n_1593);
   RAM_reg_4_74_inst : DFFX1 port map( D => n1529, CLK => n4828, Q => 
                           RAM_4_74_port, QN => n_1594);
   RAM_reg_4_73_inst : DFFX1 port map( D => n1528, CLK => n4828, Q => 
                           RAM_4_73_port, QN => n_1595);
   RAM_reg_4_72_inst : DFFX1 port map( D => n1527, CLK => n4828, Q => 
                           RAM_4_72_port, QN => n_1596);
   RAM_reg_4_71_inst : DFFX1 port map( D => n1526, CLK => n4828, Q => 
                           RAM_4_71_port, QN => n_1597);
   RAM_reg_4_70_inst : DFFX1 port map( D => n1525, CLK => n4828, Q => 
                           RAM_4_70_port, QN => n_1598);
   RAM_reg_4_69_inst : DFFX1 port map( D => n1524, CLK => n4828, Q => 
                           RAM_4_69_port, QN => n_1599);
   RAM_reg_4_68_inst : DFFX1 port map( D => n1523, CLK => n4828, Q => 
                           RAM_4_68_port, QN => n_1600);
   RAM_reg_4_67_inst : DFFX1 port map( D => n1522, CLK => n4822, Q => 
                           RAM_4_67_port, QN => n_1601);
   RAM_reg_4_66_inst : DFFX1 port map( D => n1521, CLK => n4822, Q => 
                           RAM_4_66_port, QN => n_1602);
   RAM_reg_4_65_inst : DFFX1 port map( D => n1520, CLK => n4822, Q => 
                           RAM_4_65_port, QN => n_1603);
   RAM_reg_4_64_inst : DFFX1 port map( D => n1519, CLK => n4822, Q => 
                           RAM_4_64_port, QN => n_1604);
   RAM_reg_4_63_inst : DFFX1 port map( D => n1518, CLK => n4823, Q => 
                           RAM_4_63_port, QN => n_1605);
   RAM_reg_4_62_inst : DFFX1 port map( D => n1517, CLK => n4823, Q => 
                           RAM_4_62_port, QN => n_1606);
   RAM_reg_4_61_inst : DFFX1 port map( D => n1516, CLK => n4823, Q => 
                           RAM_4_61_port, QN => n_1607);
   RAM_reg_4_60_inst : DFFX1 port map( D => n1515, CLK => n4823, Q => 
                           RAM_4_60_port, QN => n_1608);
   RAM_reg_4_59_inst : DFFX1 port map( D => n1514, CLK => n4823, Q => 
                           RAM_4_59_port, QN => n_1609);
   RAM_reg_4_58_inst : DFFX1 port map( D => n1513, CLK => n4823, Q => 
                           RAM_4_58_port, QN => n_1610);
   RAM_reg_4_57_inst : DFFX1 port map( D => n1512, CLK => n4823, Q => 
                           RAM_4_57_port, QN => n_1611);
   RAM_reg_4_56_inst : DFFX1 port map( D => n1511, CLK => n4823, Q => 
                           RAM_4_56_port, QN => n_1612);
   RAM_reg_4_55_inst : DFFX1 port map( D => n1510, CLK => n4823, Q => 
                           RAM_4_55_port, QN => n_1613);
   RAM_reg_4_54_inst : DFFX1 port map( D => n1509, CLK => n4823, Q => 
                           RAM_4_54_port, QN => n_1614);
   RAM_reg_4_53_inst : DFFX1 port map( D => n1508, CLK => n4823, Q => 
                           RAM_4_53_port, QN => n_1615);
   RAM_reg_4_52_inst : DFFX1 port map( D => n1507, CLK => n4823, Q => 
                           RAM_4_52_port, QN => n_1616);
   RAM_reg_4_51_inst : DFFX1 port map( D => n1506, CLK => n4824, Q => 
                           RAM_4_51_port, QN => n_1617);
   RAM_reg_4_50_inst : DFFX1 port map( D => n1505, CLK => n4824, Q => 
                           RAM_4_50_port, QN => n_1618);
   RAM_reg_4_49_inst : DFFX1 port map( D => n1504, CLK => n4824, Q => 
                           RAM_4_49_port, QN => n_1619);
   RAM_reg_4_48_inst : DFFX1 port map( D => n1503, CLK => n4824, Q => 
                           RAM_4_48_port, QN => n_1620);
   RAM_reg_4_47_inst : DFFX1 port map( D => n1502, CLK => n4824, Q => 
                           RAM_4_47_port, QN => n_1621);
   RAM_reg_4_46_inst : DFFX1 port map( D => n1501, CLK => n4824, Q => 
                           RAM_4_46_port, QN => n_1622);
   RAM_reg_4_45_inst : DFFX1 port map( D => n1500, CLK => n4824, Q => 
                           RAM_4_45_port, QN => n_1623);
   RAM_reg_4_44_inst : DFFX1 port map( D => n1499, CLK => n4824, Q => 
                           RAM_4_44_port, QN => n_1624);
   RAM_reg_4_43_inst : DFFX1 port map( D => n1498, CLK => n4824, Q => 
                           RAM_4_43_port, QN => n_1625);
   RAM_reg_4_42_inst : DFFX1 port map( D => n1497, CLK => n4824, Q => 
                           RAM_4_42_port, QN => n_1626);
   RAM_reg_4_41_inst : DFFX1 port map( D => n1496, CLK => n4824, Q => 
                           RAM_4_41_port, QN => n_1627);
   RAM_reg_4_40_inst : DFFX1 port map( D => n1495, CLK => n4824, Q => 
                           RAM_4_40_port, QN => n_1628);
   RAM_reg_4_39_inst : DFFX1 port map( D => n1494, CLK => n4825, Q => 
                           RAM_4_39_port, QN => n_1629);
   RAM_reg_4_38_inst : DFFX1 port map( D => n1493, CLK => n4825, Q => 
                           RAM_4_38_port, QN => n_1630);
   RAM_reg_4_37_inst : DFFX1 port map( D => n1492, CLK => n4825, Q => 
                           RAM_4_37_port, QN => n_1631);
   RAM_reg_4_36_inst : DFFX1 port map( D => n1491, CLK => n4825, Q => 
                           RAM_4_36_port, QN => n_1632);
   RAM_reg_4_35_inst : DFFX1 port map( D => n1490, CLK => n4825, Q => 
                           RAM_4_35_port, QN => n_1633);
   RAM_reg_4_34_inst : DFFX1 port map( D => n1489, CLK => n4825, Q => 
                           RAM_4_34_port, QN => n_1634);
   RAM_reg_4_33_inst : DFFX1 port map( D => n1488, CLK => n4825, Q => 
                           RAM_4_33_port, QN => n_1635);
   RAM_reg_4_32_inst : DFFX1 port map( D => n1487, CLK => n4825, Q => 
                           RAM_4_32_port, QN => n_1636);
   RAM_reg_4_31_inst : DFFX1 port map( D => n1486, CLK => n4819, Q => 
                           RAM_4_31_port, QN => n_1637);
   RAM_reg_4_30_inst : DFFX1 port map( D => n1485, CLK => n4819, Q => 
                           RAM_4_30_port, QN => n_1638);
   RAM_reg_4_29_inst : DFFX1 port map( D => n1484, CLK => n4819, Q => 
                           RAM_4_29_port, QN => n_1639);
   RAM_reg_4_28_inst : DFFX1 port map( D => n1483, CLK => n4819, Q => 
                           RAM_4_28_port, QN => n_1640);
   RAM_reg_4_27_inst : DFFX1 port map( D => n1482, CLK => n4820, Q => 
                           RAM_4_27_port, QN => n_1641);
   RAM_reg_4_26_inst : DFFX1 port map( D => n1481, CLK => n4820, Q => 
                           RAM_4_26_port, QN => n_1642);
   RAM_reg_4_25_inst : DFFX1 port map( D => n1480, CLK => n4820, Q => 
                           RAM_4_25_port, QN => n_1643);
   RAM_reg_4_24_inst : DFFX1 port map( D => n1479, CLK => n4820, Q => 
                           RAM_4_24_port, QN => n_1644);
   RAM_reg_4_23_inst : DFFX1 port map( D => n1478, CLK => n4820, Q => 
                           RAM_4_23_port, QN => n_1645);
   RAM_reg_4_22_inst : DFFX1 port map( D => n1477, CLK => n4820, Q => 
                           RAM_4_22_port, QN => n_1646);
   RAM_reg_4_21_inst : DFFX1 port map( D => n1476, CLK => n4820, Q => 
                           RAM_4_21_port, QN => n_1647);
   RAM_reg_4_20_inst : DFFX1 port map( D => n1475, CLK => n4820, Q => 
                           RAM_4_20_port, QN => n_1648);
   RAM_reg_4_19_inst : DFFX1 port map( D => n1474, CLK => n4820, Q => 
                           RAM_4_19_port, QN => n_1649);
   RAM_reg_4_18_inst : DFFX1 port map( D => n1473, CLK => n4820, Q => 
                           RAM_4_18_port, QN => n_1650);
   RAM_reg_4_17_inst : DFFX1 port map( D => n1472, CLK => n4820, Q => 
                           RAM_4_17_port, QN => n_1651);
   RAM_reg_4_16_inst : DFFX1 port map( D => n1471, CLK => n4820, Q => 
                           RAM_4_16_port, QN => n_1652);
   RAM_reg_4_15_inst : DFFX1 port map( D => n1470, CLK => n4821, Q => 
                           RAM_4_15_port, QN => n_1653);
   RAM_reg_4_14_inst : DFFX1 port map( D => n1469, CLK => n4821, Q => 
                           RAM_4_14_port, QN => n_1654);
   RAM_reg_4_13_inst : DFFX1 port map( D => n1468, CLK => n4821, Q => 
                           RAM_4_13_port, QN => n_1655);
   RAM_reg_4_12_inst : DFFX1 port map( D => n1467, CLK => n4821, Q => 
                           RAM_4_12_port, QN => n_1656);
   RAM_reg_4_11_inst : DFFX1 port map( D => n1466, CLK => n4821, Q => 
                           RAM_4_11_port, QN => n_1657);
   RAM_reg_4_10_inst : DFFX1 port map( D => n1465, CLK => n4821, Q => 
                           RAM_4_10_port, QN => n_1658);
   RAM_reg_4_9_inst : DFFX1 port map( D => n1464, CLK => n4821, Q => 
                           RAM_4_9_port, QN => n_1659);
   RAM_reg_4_8_inst : DFFX1 port map( D => n1463, CLK => n4821, Q => 
                           RAM_4_8_port, QN => n_1660);
   RAM_reg_4_7_inst : DFFX1 port map( D => n1462, CLK => n4821, Q => 
                           RAM_4_7_port, QN => n_1661);
   RAM_reg_4_6_inst : DFFX1 port map( D => n1461, CLK => n4821, Q => 
                           RAM_4_6_port, QN => n_1662);
   RAM_reg_4_5_inst : DFFX1 port map( D => n1460, CLK => n4821, Q => 
                           RAM_4_5_port, QN => n_1663);
   RAM_reg_4_4_inst : DFFX1 port map( D => n1459, CLK => n4821, Q => 
                           RAM_4_4_port, QN => n_1664);
   RAM_reg_4_3_inst : DFFX1 port map( D => n1458, CLK => n4822, Q => 
                           RAM_4_3_port, QN => n_1665);
   RAM_reg_4_2_inst : DFFX1 port map( D => n1457, CLK => n4822, Q => 
                           RAM_4_2_port, QN => n_1666);
   RAM_reg_4_1_inst : DFFX1 port map( D => n1456, CLK => n4822, Q => 
                           RAM_4_1_port, QN => n_1667);
   RAM_reg_4_0_inst : DFFX1 port map( D => n1455, CLK => n4822, Q => 
                           RAM_4_0_port, QN => n_1668);
   RAM_reg_5_127_inst : DFFX1 port map( D => n1454, CLK => n4822, Q => 
                           RAM_5_127_port, QN => n_1669);
   RAM_reg_5_126_inst : DFFX1 port map( D => n1453, CLK => n4822, Q => 
                           RAM_5_126_port, QN => n_1670);
   RAM_reg_5_125_inst : DFFX1 port map( D => n1452, CLK => n4822, Q => 
                           RAM_5_125_port, QN => n_1671);
   RAM_reg_5_124_inst : DFFX1 port map( D => n1451, CLK => n4822, Q => 
                           RAM_5_124_port, QN => n_1672);
   RAM_reg_5_123_inst : DFFX1 port map( D => n1450, CLK => n4834, Q => 
                           RAM_5_123_port, QN => n_1673);
   RAM_reg_5_122_inst : DFFX1 port map( D => n1449, CLK => n4834, Q => 
                           RAM_5_122_port, QN => n_1674);
   RAM_reg_5_121_inst : DFFX1 port map( D => n1448, CLK => n4834, Q => 
                           RAM_5_121_port, QN => n_1675);
   RAM_reg_5_120_inst : DFFX1 port map( D => n1447, CLK => n4834, Q => 
                           RAM_5_120_port, QN => n_1676);
   RAM_reg_5_119_inst : DFFX1 port map( D => n1446, CLK => n4835, Q => 
                           RAM_5_119_port, QN => n_1677);
   RAM_reg_5_118_inst : DFFX1 port map( D => n1445, CLK => n4835, Q => 
                           RAM_5_118_port, QN => n_1678);
   RAM_reg_5_117_inst : DFFX1 port map( D => n1444, CLK => n4835, Q => 
                           RAM_5_117_port, QN => n_1679);
   RAM_reg_5_116_inst : DFFX1 port map( D => n1443, CLK => n4835, Q => 
                           RAM_5_116_port, QN => n_1680);
   RAM_reg_5_115_inst : DFFX1 port map( D => n1442, CLK => n4835, Q => 
                           RAM_5_115_port, QN => n_1681);
   RAM_reg_5_114_inst : DFFX1 port map( D => n1441, CLK => n4835, Q => 
                           RAM_5_114_port, QN => n_1682);
   RAM_reg_5_113_inst : DFFX1 port map( D => n1440, CLK => n4835, Q => 
                           RAM_5_113_port, QN => n_1683);
   RAM_reg_5_112_inst : DFFX1 port map( D => n1439, CLK => n4835, Q => 
                           RAM_5_112_port, QN => n_1684);
   RAM_reg_5_111_inst : DFFX1 port map( D => n1438, CLK => n4835, Q => 
                           RAM_5_111_port, QN => n_1685);
   RAM_reg_5_110_inst : DFFX1 port map( D => n1437, CLK => n4835, Q => 
                           RAM_5_110_port, QN => n_1686);
   RAM_reg_5_109_inst : DFFX1 port map( D => n1436, CLK => n4835, Q => 
                           RAM_5_109_port, QN => n_1687);
   RAM_reg_5_108_inst : DFFX1 port map( D => n1435, CLK => n4835, Q => 
                           RAM_5_108_port, QN => n_1688);
   RAM_reg_5_107_inst : DFFX1 port map( D => n1434, CLK => n4836, Q => 
                           RAM_5_107_port, QN => n_1689);
   RAM_reg_5_106_inst : DFFX1 port map( D => n1433, CLK => n4836, Q => 
                           RAM_5_106_port, QN => n_1690);
   RAM_reg_5_105_inst : DFFX1 port map( D => n1432, CLK => n4836, Q => 
                           RAM_5_105_port, QN => n_1691);
   RAM_reg_5_104_inst : DFFX1 port map( D => n1431, CLK => n4836, Q => 
                           RAM_5_104_port, QN => n_1692);
   RAM_reg_5_103_inst : DFFX1 port map( D => n1430, CLK => n4836, Q => 
                           RAM_5_103_port, QN => n_1693);
   RAM_reg_5_102_inst : DFFX1 port map( D => n1429, CLK => n4836, Q => 
                           RAM_5_102_port, QN => n_1694);
   RAM_reg_5_101_inst : DFFX1 port map( D => n1428, CLK => n4836, Q => 
                           RAM_5_101_port, QN => n_1695);
   RAM_reg_5_100_inst : DFFX1 port map( D => n1427, CLK => n4836, Q => 
                           RAM_5_100_port, QN => n_1696);
   RAM_reg_5_99_inst : DFFX1 port map( D => n1426, CLK => n4836, Q => 
                           RAM_5_99_port, QN => n_1697);
   RAM_reg_5_98_inst : DFFX1 port map( D => n1425, CLK => n4836, Q => 
                           RAM_5_98_port, QN => n_1698);
   RAM_reg_5_97_inst : DFFX1 port map( D => n1424, CLK => n4836, Q => 
                           RAM_5_97_port, QN => n_1699);
   RAM_reg_5_96_inst : DFFX1 port map( D => n1423, CLK => n4836, Q => 
                           RAM_5_96_port, QN => n_1700);
   RAM_reg_5_95_inst : DFFX1 port map( D => n1422, CLK => n4837, Q => 
                           RAM_5_95_port, QN => n_1701);
   RAM_reg_5_94_inst : DFFX1 port map( D => n1421, CLK => n4837, Q => 
                           RAM_5_94_port, QN => n_1702);
   RAM_reg_5_93_inst : DFFX1 port map( D => n1420, CLK => n4837, Q => 
                           RAM_5_93_port, QN => n_1703);
   RAM_reg_5_92_inst : DFFX1 port map( D => n1419, CLK => n4837, Q => 
                           RAM_5_92_port, QN => n_1704);
   RAM_reg_5_91_inst : DFFX1 port map( D => n1418, CLK => n4837, Q => 
                           RAM_5_91_port, QN => n_1705);
   RAM_reg_5_90_inst : DFFX1 port map( D => n1417, CLK => n4837, Q => 
                           RAM_5_90_port, QN => n_1706);
   RAM_reg_5_89_inst : DFFX1 port map( D => n1416, CLK => n4837, Q => 
                           RAM_5_89_port, QN => n_1707);
   RAM_reg_5_88_inst : DFFX1 port map( D => n1415, CLK => n4837, Q => 
                           RAM_5_88_port, QN => n_1708);
   RAM_reg_5_87_inst : DFFX1 port map( D => n1414, CLK => n4831, Q => 
                           RAM_5_87_port, QN => n_1709);
   RAM_reg_5_86_inst : DFFX1 port map( D => n1413, CLK => n4831, Q => 
                           RAM_5_86_port, QN => n_1710);
   RAM_reg_5_85_inst : DFFX1 port map( D => n1412, CLK => n4831, Q => 
                           RAM_5_85_port, QN => n_1711);
   RAM_reg_5_84_inst : DFFX1 port map( D => n1411, CLK => n4831, Q => 
                           RAM_5_84_port, QN => n_1712);
   RAM_reg_5_83_inst : DFFX1 port map( D => n1410, CLK => n4832, Q => 
                           RAM_5_83_port, QN => n_1713);
   RAM_reg_5_82_inst : DFFX1 port map( D => n1409, CLK => n4832, Q => 
                           RAM_5_82_port, QN => n_1714);
   RAM_reg_5_81_inst : DFFX1 port map( D => n1408, CLK => n4832, Q => 
                           RAM_5_81_port, QN => n_1715);
   RAM_reg_5_80_inst : DFFX1 port map( D => n1407, CLK => n4832, Q => 
                           RAM_5_80_port, QN => n_1716);
   RAM_reg_5_79_inst : DFFX1 port map( D => n1406, CLK => n4832, Q => 
                           RAM_5_79_port, QN => n_1717);
   RAM_reg_5_78_inst : DFFX1 port map( D => n1405, CLK => n4832, Q => 
                           RAM_5_78_port, QN => n_1718);
   RAM_reg_5_77_inst : DFFX1 port map( D => n1404, CLK => n4832, Q => 
                           RAM_5_77_port, QN => n_1719);
   RAM_reg_5_76_inst : DFFX1 port map( D => n1403, CLK => n4832, Q => 
                           RAM_5_76_port, QN => n_1720);
   RAM_reg_5_75_inst : DFFX1 port map( D => n1402, CLK => n4832, Q => 
                           RAM_5_75_port, QN => n_1721);
   RAM_reg_5_74_inst : DFFX1 port map( D => n1401, CLK => n4832, Q => 
                           RAM_5_74_port, QN => n_1722);
   RAM_reg_5_73_inst : DFFX1 port map( D => n1400, CLK => n4832, Q => 
                           RAM_5_73_port, QN => n_1723);
   RAM_reg_5_72_inst : DFFX1 port map( D => n1399, CLK => n4832, Q => 
                           RAM_5_72_port, QN => n_1724);
   RAM_reg_5_71_inst : DFFX1 port map( D => n1398, CLK => n4833, Q => 
                           RAM_5_71_port, QN => n_1725);
   RAM_reg_5_70_inst : DFFX1 port map( D => n1397, CLK => n4833, Q => 
                           RAM_5_70_port, QN => n_1726);
   RAM_reg_5_69_inst : DFFX1 port map( D => n1396, CLK => n4833, Q => 
                           RAM_5_69_port, QN => n_1727);
   RAM_reg_5_68_inst : DFFX1 port map( D => n1395, CLK => n4833, Q => 
                           RAM_5_68_port, QN => n_1728);
   RAM_reg_5_67_inst : DFFX1 port map( D => n1394, CLK => n4833, Q => 
                           RAM_5_67_port, QN => n_1729);
   RAM_reg_5_66_inst : DFFX1 port map( D => n1393, CLK => n4833, Q => 
                           RAM_5_66_port, QN => n_1730);
   RAM_reg_5_65_inst : DFFX1 port map( D => n1392, CLK => n4833, Q => 
                           RAM_5_65_port, QN => n_1731);
   RAM_reg_5_64_inst : DFFX1 port map( D => n1391, CLK => n4833, Q => 
                           RAM_5_64_port, QN => n_1732);
   RAM_reg_5_63_inst : DFFX1 port map( D => n1390, CLK => n4833, Q => 
                           RAM_5_63_port, QN => n_1733);
   RAM_reg_5_62_inst : DFFX1 port map( D => n1389, CLK => n4833, Q => 
                           RAM_5_62_port, QN => n_1734);
   RAM_reg_5_61_inst : DFFX1 port map( D => n1388, CLK => n4833, Q => 
                           RAM_5_61_port, QN => n_1735);
   RAM_reg_5_60_inst : DFFX1 port map( D => n1387, CLK => n4833, Q => 
                           RAM_5_60_port, QN => n_1736);
   RAM_reg_5_59_inst : DFFX1 port map( D => n1386, CLK => n4834, Q => 
                           RAM_5_59_port, QN => n_1737);
   RAM_reg_5_58_inst : DFFX1 port map( D => n1385, CLK => n4834, Q => 
                           RAM_5_58_port, QN => n_1738);
   RAM_reg_5_57_inst : DFFX1 port map( D => n1384, CLK => n4834, Q => 
                           RAM_5_57_port, QN => n_1739);
   RAM_reg_5_56_inst : DFFX1 port map( D => n1383, CLK => n4834, Q => 
                           RAM_5_56_port, QN => n_1740);
   RAM_reg_5_55_inst : DFFX1 port map( D => n1382, CLK => n4834, Q => 
                           RAM_5_55_port, QN => n_1741);
   RAM_reg_5_54_inst : DFFX1 port map( D => n1381, CLK => n4834, Q => 
                           RAM_5_54_port, QN => n_1742);
   RAM_reg_5_53_inst : DFFX1 port map( D => n1380, CLK => n4834, Q => 
                           RAM_5_53_port, QN => n_1743);
   RAM_reg_5_52_inst : DFFX1 port map( D => n1379, CLK => n4834, Q => 
                           RAM_5_52_port, QN => n_1744);
   RAM_reg_5_51_inst : DFFX1 port map( D => n1378, CLK => n4828, Q => 
                           RAM_5_51_port, QN => n_1745);
   RAM_reg_5_50_inst : DFFX1 port map( D => n1377, CLK => n4828, Q => 
                           RAM_5_50_port, QN => n_1746);
   RAM_reg_5_49_inst : DFFX1 port map( D => n1376, CLK => n4828, Q => 
                           RAM_5_49_port, QN => n_1747);
   RAM_reg_5_48_inst : DFFX1 port map( D => n1375, CLK => n4828, Q => 
                           RAM_5_48_port, QN => n_1748);
   RAM_reg_5_47_inst : DFFX1 port map( D => n1374, CLK => n4829, Q => 
                           RAM_5_47_port, QN => n_1749);
   RAM_reg_5_46_inst : DFFX1 port map( D => n1373, CLK => n4829, Q => 
                           RAM_5_46_port, QN => n_1750);
   RAM_reg_5_45_inst : DFFX1 port map( D => n1372, CLK => n4829, Q => 
                           RAM_5_45_port, QN => n_1751);
   RAM_reg_5_44_inst : DFFX1 port map( D => n1371, CLK => n4829, Q => 
                           RAM_5_44_port, QN => n_1752);
   RAM_reg_5_43_inst : DFFX1 port map( D => n1370, CLK => n4829, Q => 
                           RAM_5_43_port, QN => n_1753);
   RAM_reg_5_42_inst : DFFX1 port map( D => n1369, CLK => n4829, Q => 
                           RAM_5_42_port, QN => n_1754);
   RAM_reg_5_41_inst : DFFX1 port map( D => n1368, CLK => n4829, Q => 
                           RAM_5_41_port, QN => n_1755);
   RAM_reg_5_40_inst : DFFX1 port map( D => n1367, CLK => n4829, Q => 
                           RAM_5_40_port, QN => n_1756);
   RAM_reg_5_39_inst : DFFX1 port map( D => n1366, CLK => n4829, Q => 
                           RAM_5_39_port, QN => n_1757);
   RAM_reg_5_38_inst : DFFX1 port map( D => n1365, CLK => n4829, Q => 
                           RAM_5_38_port, QN => n_1758);
   RAM_reg_5_37_inst : DFFX1 port map( D => n1364, CLK => n4829, Q => 
                           RAM_5_37_port, QN => n_1759);
   RAM_reg_5_36_inst : DFFX1 port map( D => n1363, CLK => n4829, Q => 
                           RAM_5_36_port, QN => n_1760);
   RAM_reg_5_35_inst : DFFX1 port map( D => n1362, CLK => n4830, Q => 
                           RAM_5_35_port, QN => n_1761);
   RAM_reg_5_34_inst : DFFX1 port map( D => n1361, CLK => n4830, Q => 
                           RAM_5_34_port, QN => n_1762);
   RAM_reg_5_33_inst : DFFX1 port map( D => n1360, CLK => n4830, Q => 
                           RAM_5_33_port, QN => n_1763);
   RAM_reg_5_32_inst : DFFX1 port map( D => n1359, CLK => n4830, Q => 
                           RAM_5_32_port, QN => n_1764);
   RAM_reg_5_31_inst : DFFX1 port map( D => n1358, CLK => n4830, Q => 
                           RAM_5_31_port, QN => n_1765);
   RAM_reg_5_30_inst : DFFX1 port map( D => n1357, CLK => n4830, Q => 
                           RAM_5_30_port, QN => n_1766);
   RAM_reg_5_29_inst : DFFX1 port map( D => n1356, CLK => n4830, Q => 
                           RAM_5_29_port, QN => n_1767);
   RAM_reg_5_28_inst : DFFX1 port map( D => n1355, CLK => n4830, Q => 
                           RAM_5_28_port, QN => n_1768);
   RAM_reg_5_27_inst : DFFX1 port map( D => n1354, CLK => n4830, Q => 
                           RAM_5_27_port, QN => n_1769);
   RAM_reg_5_26_inst : DFFX1 port map( D => n1353, CLK => n4830, Q => 
                           RAM_5_26_port, QN => n_1770);
   RAM_reg_5_25_inst : DFFX1 port map( D => n1352, CLK => n4830, Q => 
                           RAM_5_25_port, QN => n_1771);
   RAM_reg_5_24_inst : DFFX1 port map( D => n1351, CLK => n4830, Q => 
                           RAM_5_24_port, QN => n_1772);
   RAM_reg_5_23_inst : DFFX1 port map( D => n1350, CLK => n4831, Q => 
                           RAM_5_23_port, QN => n_1773);
   RAM_reg_5_22_inst : DFFX1 port map( D => n1349, CLK => n4831, Q => 
                           RAM_5_22_port, QN => n_1774);
   RAM_reg_5_21_inst : DFFX1 port map( D => n1348, CLK => n4831, Q => 
                           RAM_5_21_port, QN => n_1775);
   RAM_reg_5_20_inst : DFFX1 port map( D => n1347, CLK => n4831, Q => 
                           RAM_5_20_port, QN => n_1776);
   RAM_reg_5_19_inst : DFFX1 port map( D => n1346, CLK => n4831, Q => 
                           RAM_5_19_port, QN => n_1777);
   RAM_reg_5_18_inst : DFFX1 port map( D => n1345, CLK => n4831, Q => 
                           RAM_5_18_port, QN => n_1778);
   RAM_reg_5_17_inst : DFFX1 port map( D => n1344, CLK => n4831, Q => 
                           RAM_5_17_port, QN => n_1779);
   RAM_reg_5_16_inst : DFFX1 port map( D => n1343, CLK => n4831, Q => 
                           RAM_5_16_port, QN => n_1780);
   RAM_reg_5_15_inst : DFFX1 port map( D => n1342, CLK => n4843, Q => 
                           RAM_5_15_port, QN => n_1781);
   RAM_reg_5_14_inst : DFFX1 port map( D => n1341, CLK => n4843, Q => 
                           RAM_5_14_port, QN => n_1782);
   RAM_reg_5_13_inst : DFFX1 port map( D => n1340, CLK => n4843, Q => 
                           RAM_5_13_port, QN => n_1783);
   RAM_reg_5_12_inst : DFFX1 port map( D => n1339, CLK => n4843, Q => 
                           RAM_5_12_port, QN => n_1784);
   RAM_reg_5_11_inst : DFFX1 port map( D => n1338, CLK => n4844, Q => 
                           RAM_5_11_port, QN => n_1785);
   RAM_reg_5_10_inst : DFFX1 port map( D => n1337, CLK => n4844, Q => 
                           RAM_5_10_port, QN => n_1786);
   RAM_reg_5_9_inst : DFFX1 port map( D => n1336, CLK => n4844, Q => 
                           RAM_5_9_port, QN => n_1787);
   RAM_reg_5_8_inst : DFFX1 port map( D => n1335, CLK => n4844, Q => 
                           RAM_5_8_port, QN => n_1788);
   RAM_reg_5_7_inst : DFFX1 port map( D => n1334, CLK => n4844, Q => 
                           RAM_5_7_port, QN => n_1789);
   RAM_reg_5_6_inst : DFFX1 port map( D => n1333, CLK => n4844, Q => 
                           RAM_5_6_port, QN => n_1790);
   RAM_reg_5_5_inst : DFFX1 port map( D => n1332, CLK => n4844, Q => 
                           RAM_5_5_port, QN => n_1791);
   RAM_reg_5_4_inst : DFFX1 port map( D => n1331, CLK => n4844, Q => 
                           RAM_5_4_port, QN => n_1792);
   RAM_reg_5_3_inst : DFFX1 port map( D => n1330, CLK => n4844, Q => 
                           RAM_5_3_port, QN => n_1793);
   RAM_reg_5_2_inst : DFFX1 port map( D => n1329, CLK => n4844, Q => 
                           RAM_5_2_port, QN => n_1794);
   RAM_reg_5_1_inst : DFFX1 port map( D => n1328, CLK => n4844, Q => 
                           RAM_5_1_port, QN => n_1795);
   RAM_reg_5_0_inst : DFFX1 port map( D => n1327, CLK => n4844, Q => 
                           RAM_5_0_port, QN => n_1796);
   RAM_reg_6_127_inst : DFFX1 port map( D => n1326, CLK => n4845, Q => 
                           RAM_6_127_port, QN => n_1797);
   RAM_reg_6_126_inst : DFFX1 port map( D => n1325, CLK => n4845, Q => 
                           RAM_6_126_port, QN => n_1798);
   RAM_reg_6_125_inst : DFFX1 port map( D => n1324, CLK => n4845, Q => 
                           RAM_6_125_port, QN => n_1799);
   RAM_reg_6_124_inst : DFFX1 port map( D => n1323, CLK => n4845, Q => 
                           RAM_6_124_port, QN => n_1800);
   RAM_reg_6_123_inst : DFFX1 port map( D => n1322, CLK => n4845, Q => 
                           RAM_6_123_port, QN => n_1801);
   RAM_reg_6_122_inst : DFFX1 port map( D => n1321, CLK => n4845, Q => 
                           RAM_6_122_port, QN => n_1802);
   RAM_reg_6_121_inst : DFFX1 port map( D => n1320, CLK => n4845, Q => 
                           RAM_6_121_port, QN => n_1803);
   RAM_reg_6_120_inst : DFFX1 port map( D => n1319, CLK => n4845, Q => 
                           RAM_6_120_port, QN => n_1804);
   RAM_reg_6_119_inst : DFFX1 port map( D => n1318, CLK => n4845, Q => 
                           RAM_6_119_port, QN => n_1805);
   RAM_reg_6_118_inst : DFFX1 port map( D => n1317, CLK => n4845, Q => 
                           RAM_6_118_port, QN => n_1806);
   RAM_reg_6_117_inst : DFFX1 port map( D => n1316, CLK => n4845, Q => 
                           RAM_6_117_port, QN => n_1807);
   RAM_reg_6_116_inst : DFFX1 port map( D => n1315, CLK => n4845, Q => 
                           RAM_6_116_port, QN => n_1808);
   RAM_reg_6_115_inst : DFFX1 port map( D => n1314, CLK => n4846, Q => 
                           RAM_6_115_port, QN => n_1809);
   RAM_reg_6_114_inst : DFFX1 port map( D => n1313, CLK => n4846, Q => 
                           RAM_6_114_port, QN => n_1810);
   RAM_reg_6_113_inst : DFFX1 port map( D => n1312, CLK => n4846, Q => 
                           RAM_6_113_port, QN => n_1811);
   RAM_reg_6_112_inst : DFFX1 port map( D => n1311, CLK => n4846, Q => 
                           RAM_6_112_port, QN => n_1812);
   RAM_reg_6_111_inst : DFFX1 port map( D => n1310, CLK => n4846, Q => 
                           RAM_6_111_port, QN => n_1813);
   RAM_reg_6_110_inst : DFFX1 port map( D => n1309, CLK => n4846, Q => 
                           RAM_6_110_port, QN => n_1814);
   RAM_reg_6_109_inst : DFFX1 port map( D => n1308, CLK => n4846, Q => 
                           RAM_6_109_port, QN => n_1815);
   RAM_reg_6_108_inst : DFFX1 port map( D => n1307, CLK => n4846, Q => 
                           RAM_6_108_port, QN => n_1816);
   RAM_reg_6_107_inst : DFFX1 port map( D => n1306, CLK => n4840, Q => 
                           RAM_6_107_port, QN => n_1817);
   RAM_reg_6_106_inst : DFFX1 port map( D => n1305, CLK => n4840, Q => 
                           RAM_6_106_port, QN => n_1818);
   RAM_reg_6_105_inst : DFFX1 port map( D => n1304, CLK => n4840, Q => 
                           RAM_6_105_port, QN => n_1819);
   RAM_reg_6_104_inst : DFFX1 port map( D => n1303, CLK => n4840, Q => 
                           RAM_6_104_port, QN => n_1820);
   RAM_reg_6_103_inst : DFFX1 port map( D => n1302, CLK => n4841, Q => 
                           RAM_6_103_port, QN => n_1821);
   RAM_reg_6_102_inst : DFFX1 port map( D => n1301, CLK => n4841, Q => 
                           RAM_6_102_port, QN => n_1822);
   RAM_reg_6_101_inst : DFFX1 port map( D => n1300, CLK => n4841, Q => 
                           RAM_6_101_port, QN => n_1823);
   RAM_reg_6_100_inst : DFFX1 port map( D => n1299, CLK => n4841, Q => 
                           RAM_6_100_port, QN => n_1824);
   RAM_reg_6_99_inst : DFFX1 port map( D => n1298, CLK => n4841, Q => 
                           RAM_6_99_port, QN => n_1825);
   RAM_reg_6_98_inst : DFFX1 port map( D => n1297, CLK => n4841, Q => 
                           RAM_6_98_port, QN => n_1826);
   RAM_reg_6_97_inst : DFFX1 port map( D => n1296, CLK => n4841, Q => 
                           RAM_6_97_port, QN => n_1827);
   RAM_reg_6_96_inst : DFFX1 port map( D => n1295, CLK => n4841, Q => 
                           RAM_6_96_port, QN => n_1828);
   RAM_reg_6_95_inst : DFFX1 port map( D => n1294, CLK => n4841, Q => 
                           RAM_6_95_port, QN => n_1829);
   RAM_reg_6_94_inst : DFFX1 port map( D => n1293, CLK => n4841, Q => 
                           RAM_6_94_port, QN => n_1830);
   RAM_reg_6_93_inst : DFFX1 port map( D => n1292, CLK => n4841, Q => 
                           RAM_6_93_port, QN => n_1831);
   RAM_reg_6_92_inst : DFFX1 port map( D => n1291, CLK => n4841, Q => 
                           RAM_6_92_port, QN => n_1832);
   RAM_reg_6_91_inst : DFFX1 port map( D => n1290, CLK => n4842, Q => 
                           RAM_6_91_port, QN => n_1833);
   RAM_reg_6_90_inst : DFFX1 port map( D => n1289, CLK => n4842, Q => 
                           RAM_6_90_port, QN => n_1834);
   RAM_reg_6_89_inst : DFFX1 port map( D => n1288, CLK => n4842, Q => 
                           RAM_6_89_port, QN => n_1835);
   RAM_reg_6_88_inst : DFFX1 port map( D => n1287, CLK => n4842, Q => 
                           RAM_6_88_port, QN => n_1836);
   RAM_reg_6_87_inst : DFFX1 port map( D => n1286, CLK => n4842, Q => 
                           RAM_6_87_port, QN => n_1837);
   RAM_reg_6_86_inst : DFFX1 port map( D => n1285, CLK => n4842, Q => 
                           RAM_6_86_port, QN => n_1838);
   RAM_reg_6_85_inst : DFFX1 port map( D => n1284, CLK => n4842, Q => 
                           RAM_6_85_port, QN => n_1839);
   RAM_reg_6_84_inst : DFFX1 port map( D => n1283, CLK => n4842, Q => 
                           RAM_6_84_port, QN => n_1840);
   RAM_reg_6_83_inst : DFFX1 port map( D => n1282, CLK => n4842, Q => 
                           RAM_6_83_port, QN => n_1841);
   RAM_reg_6_82_inst : DFFX1 port map( D => n1281, CLK => n4842, Q => 
                           RAM_6_82_port, QN => n_1842);
   RAM_reg_6_81_inst : DFFX1 port map( D => n1280, CLK => n4842, Q => 
                           RAM_6_81_port, QN => n_1843);
   RAM_reg_6_80_inst : DFFX1 port map( D => n1279, CLK => n4842, Q => 
                           RAM_6_80_port, QN => n_1844);
   RAM_reg_6_79_inst : DFFX1 port map( D => n1278, CLK => n4843, Q => 
                           RAM_6_79_port, QN => n_1845);
   RAM_reg_6_78_inst : DFFX1 port map( D => n1277, CLK => n4843, Q => 
                           RAM_6_78_port, QN => n_1846);
   RAM_reg_6_77_inst : DFFX1 port map( D => n1276, CLK => n4843, Q => 
                           RAM_6_77_port, QN => n_1847);
   RAM_reg_6_76_inst : DFFX1 port map( D => n1275, CLK => n4843, Q => 
                           RAM_6_76_port, QN => n_1848);
   RAM_reg_6_75_inst : DFFX1 port map( D => n1274, CLK => n4843, Q => 
                           RAM_6_75_port, QN => n_1849);
   RAM_reg_6_74_inst : DFFX1 port map( D => n1273, CLK => n4843, Q => 
                           RAM_6_74_port, QN => n_1850);
   RAM_reg_6_73_inst : DFFX1 port map( D => n1272, CLK => n4843, Q => 
                           RAM_6_73_port, QN => n_1851);
   RAM_reg_6_72_inst : DFFX1 port map( D => n1271, CLK => n4843, Q => 
                           RAM_6_72_port, QN => n_1852);
   RAM_reg_6_71_inst : DFFX1 port map( D => n1270, CLK => n4837, Q => 
                           RAM_6_71_port, QN => n_1853);
   RAM_reg_6_70_inst : DFFX1 port map( D => n1269, CLK => n4837, Q => 
                           RAM_6_70_port, QN => n_1854);
   RAM_reg_6_69_inst : DFFX1 port map( D => n1268, CLK => n4837, Q => 
                           RAM_6_69_port, QN => n_1855);
   RAM_reg_6_68_inst : DFFX1 port map( D => n1267, CLK => n4837, Q => 
                           RAM_6_68_port, QN => n_1856);
   RAM_reg_6_67_inst : DFFX1 port map( D => n1266, CLK => n4838, Q => 
                           RAM_6_67_port, QN => n_1857);
   RAM_reg_6_66_inst : DFFX1 port map( D => n1265, CLK => n4838, Q => 
                           RAM_6_66_port, QN => n_1858);
   RAM_reg_6_65_inst : DFFX1 port map( D => n1264, CLK => n4838, Q => 
                           RAM_6_65_port, QN => n_1859);
   RAM_reg_6_64_inst : DFFX1 port map( D => n1263, CLK => n4838, Q => 
                           RAM_6_64_port, QN => n_1860);
   RAM_reg_6_63_inst : DFFX1 port map( D => n1262, CLK => n4838, Q => 
                           RAM_6_63_port, QN => n_1861);
   RAM_reg_6_62_inst : DFFX1 port map( D => n1261, CLK => n4838, Q => 
                           RAM_6_62_port, QN => n_1862);
   RAM_reg_6_61_inst : DFFX1 port map( D => n1260, CLK => n4838, Q => 
                           RAM_6_61_port, QN => n_1863);
   RAM_reg_6_60_inst : DFFX1 port map( D => n1259, CLK => n4838, Q => 
                           RAM_6_60_port, QN => n_1864);
   RAM_reg_6_59_inst : DFFX1 port map( D => n1258, CLK => n4838, Q => 
                           RAM_6_59_port, QN => n_1865);
   RAM_reg_6_58_inst : DFFX1 port map( D => n1257, CLK => n4838, Q => 
                           RAM_6_58_port, QN => n_1866);
   RAM_reg_6_57_inst : DFFX1 port map( D => n1256, CLK => n4838, Q => 
                           RAM_6_57_port, QN => n_1867);
   RAM_reg_6_56_inst : DFFX1 port map( D => n1255, CLK => n4838, Q => 
                           RAM_6_56_port, QN => n_1868);
   RAM_reg_6_55_inst : DFFX1 port map( D => n1254, CLK => n4839, Q => 
                           RAM_6_55_port, QN => n_1869);
   RAM_reg_6_54_inst : DFFX1 port map( D => n1253, CLK => n4839, Q => 
                           RAM_6_54_port, QN => n_1870);
   RAM_reg_6_53_inst : DFFX1 port map( D => n1252, CLK => n4839, Q => 
                           RAM_6_53_port, QN => n_1871);
   RAM_reg_6_52_inst : DFFX1 port map( D => n1251, CLK => n4839, Q => 
                           RAM_6_52_port, QN => n_1872);
   RAM_reg_6_51_inst : DFFX1 port map( D => n1250, CLK => n4839, Q => 
                           RAM_6_51_port, QN => n_1873);
   RAM_reg_6_50_inst : DFFX1 port map( D => n1249, CLK => n4839, Q => 
                           RAM_6_50_port, QN => n_1874);
   RAM_reg_6_49_inst : DFFX1 port map( D => n1248, CLK => n4839, Q => 
                           RAM_6_49_port, QN => n_1875);
   RAM_reg_6_48_inst : DFFX1 port map( D => n1247, CLK => n4839, Q => 
                           RAM_6_48_port, QN => n_1876);
   RAM_reg_6_47_inst : DFFX1 port map( D => n1246, CLK => n4839, Q => 
                           RAM_6_47_port, QN => n_1877);
   RAM_reg_6_46_inst : DFFX1 port map( D => n1245, CLK => n4839, Q => 
                           RAM_6_46_port, QN => n_1878);
   RAM_reg_6_45_inst : DFFX1 port map( D => n1244, CLK => n4839, Q => 
                           RAM_6_45_port, QN => n_1879);
   RAM_reg_6_44_inst : DFFX1 port map( D => n1243, CLK => n4839, Q => 
                           RAM_6_44_port, QN => n_1880);
   RAM_reg_6_43_inst : DFFX1 port map( D => n1242, CLK => n4840, Q => 
                           RAM_6_43_port, QN => n_1881);
   RAM_reg_6_42_inst : DFFX1 port map( D => n1241, CLK => n4840, Q => 
                           RAM_6_42_port, QN => n_1882);
   RAM_reg_6_41_inst : DFFX1 port map( D => n1240, CLK => n4840, Q => 
                           RAM_6_41_port, QN => n_1883);
   RAM_reg_6_40_inst : DFFX1 port map( D => n1239, CLK => n4840, Q => 
                           RAM_6_40_port, QN => n_1884);
   RAM_reg_6_39_inst : DFFX1 port map( D => n1238, CLK => n4840, Q => 
                           RAM_6_39_port, QN => n_1885);
   RAM_reg_6_38_inst : DFFX1 port map( D => n1237, CLK => n4840, Q => 
                           RAM_6_38_port, QN => n_1886);
   RAM_reg_6_37_inst : DFFX1 port map( D => n1236, CLK => n4840, Q => 
                           RAM_6_37_port, QN => n_1887);
   RAM_reg_6_36_inst : DFFX1 port map( D => n1235, CLK => n4840, Q => 
                           RAM_6_36_port, QN => n_1888);
   RAM_reg_6_35_inst : DFFX1 port map( D => n1234, CLK => n4852, Q => 
                           RAM_6_35_port, QN => n_1889);
   RAM_reg_6_34_inst : DFFX1 port map( D => n1233, CLK => n4852, Q => 
                           RAM_6_34_port, QN => n_1890);
   RAM_reg_6_33_inst : DFFX1 port map( D => n1232, CLK => n4852, Q => 
                           RAM_6_33_port, QN => n_1891);
   RAM_reg_6_32_inst : DFFX1 port map( D => n1231, CLK => n4852, Q => 
                           RAM_6_32_port, QN => n_1892);
   RAM_reg_6_31_inst : DFFX1 port map( D => n1230, CLK => n4853, Q => 
                           RAM_6_31_port, QN => n_1893);
   RAM_reg_6_30_inst : DFFX1 port map( D => n1229, CLK => n4853, Q => 
                           RAM_6_30_port, QN => n_1894);
   RAM_reg_6_29_inst : DFFX1 port map( D => n1228, CLK => n4853, Q => 
                           RAM_6_29_port, QN => n_1895);
   RAM_reg_6_28_inst : DFFX1 port map( D => n1227, CLK => n4853, Q => 
                           RAM_6_28_port, QN => n_1896);
   RAM_reg_6_27_inst : DFFX1 port map( D => n1226, CLK => n4853, Q => 
                           RAM_6_27_port, QN => n_1897);
   RAM_reg_6_26_inst : DFFX1 port map( D => n1225, CLK => n4853, Q => 
                           RAM_6_26_port, QN => n_1898);
   RAM_reg_6_25_inst : DFFX1 port map( D => n1224, CLK => n4853, Q => 
                           RAM_6_25_port, QN => n_1899);
   RAM_reg_6_24_inst : DFFX1 port map( D => n1223, CLK => n4853, Q => 
                           RAM_6_24_port, QN => n_1900);
   RAM_reg_6_23_inst : DFFX1 port map( D => n1222, CLK => n4853, Q => 
                           RAM_6_23_port, QN => n_1901);
   RAM_reg_6_22_inst : DFFX1 port map( D => n1221, CLK => n4853, Q => 
                           RAM_6_22_port, QN => n_1902);
   RAM_reg_6_21_inst : DFFX1 port map( D => n1220, CLK => n4853, Q => 
                           RAM_6_21_port, QN => n_1903);
   RAM_reg_6_20_inst : DFFX1 port map( D => n1219, CLK => n4853, Q => 
                           RAM_6_20_port, QN => n_1904);
   RAM_reg_6_19_inst : DFFX1 port map( D => n1218, CLK => n4854, Q => 
                           RAM_6_19_port, QN => n_1905);
   RAM_reg_6_18_inst : DFFX1 port map( D => n1217, CLK => n4854, Q => 
                           RAM_6_18_port, QN => n_1906);
   RAM_reg_6_17_inst : DFFX1 port map( D => n1216, CLK => n4854, Q => 
                           RAM_6_17_port, QN => n_1907);
   RAM_reg_6_16_inst : DFFX1 port map( D => n1215, CLK => n4854, Q => 
                           RAM_6_16_port, QN => n_1908);
   RAM_reg_6_15_inst : DFFX1 port map( D => n1214, CLK => n4854, Q => 
                           RAM_6_15_port, QN => n_1909);
   RAM_reg_6_14_inst : DFFX1 port map( D => n1213, CLK => n4854, Q => 
                           RAM_6_14_port, QN => n_1910);
   RAM_reg_6_13_inst : DFFX1 port map( D => n1212, CLK => n4854, Q => 
                           RAM_6_13_port, QN => n_1911);
   RAM_reg_6_12_inst : DFFX1 port map( D => n1211, CLK => n4854, Q => 
                           RAM_6_12_port, QN => n_1912);
   RAM_reg_6_11_inst : DFFX1 port map( D => n1210, CLK => n4854, Q => 
                           RAM_6_11_port, QN => n_1913);
   RAM_reg_6_10_inst : DFFX1 port map( D => n1209, CLK => n4854, Q => 
                           RAM_6_10_port, QN => n_1914);
   RAM_reg_6_9_inst : DFFX1 port map( D => n1208, CLK => n4854, Q => 
                           RAM_6_9_port, QN => n_1915);
   RAM_reg_6_8_inst : DFFX1 port map( D => n1207, CLK => n4854, Q => 
                           RAM_6_8_port, QN => n_1916);
   RAM_reg_6_7_inst : DFFX1 port map( D => n1206, CLK => n4855, Q => 
                           RAM_6_7_port, QN => n_1917);
   RAM_reg_6_6_inst : DFFX1 port map( D => n1205, CLK => n4855, Q => 
                           RAM_6_6_port, QN => n_1918);
   RAM_reg_6_5_inst : DFFX1 port map( D => n1204, CLK => n4855, Q => 
                           RAM_6_5_port, QN => n_1919);
   RAM_reg_6_4_inst : DFFX1 port map( D => n1203, CLK => n4855, Q => 
                           RAM_6_4_port, QN => n_1920);
   RAM_reg_6_3_inst : DFFX1 port map( D => n1202, CLK => n4855, Q => 
                           RAM_6_3_port, QN => n_1921);
   RAM_reg_6_2_inst : DFFX1 port map( D => n1201, CLK => n4855, Q => 
                           RAM_6_2_port, QN => n_1922);
   RAM_reg_6_1_inst : DFFX1 port map( D => n1200, CLK => n4855, Q => 
                           RAM_6_1_port, QN => n_1923);
   RAM_reg_6_0_inst : DFFX1 port map( D => n1199, CLK => n4855, Q => 
                           RAM_6_0_port, QN => n_1924);
   RAM_reg_7_127_inst : DFFX1 port map( D => n1198, CLK => n4849, Q => 
                           RAM_7_127_port, QN => n_1925);
   RAM_reg_7_126_inst : DFFX1 port map( D => n1197, CLK => n4849, Q => 
                           RAM_7_126_port, QN => n_1926);
   RAM_reg_7_125_inst : DFFX1 port map( D => n1196, CLK => n4849, Q => 
                           RAM_7_125_port, QN => n_1927);
   RAM_reg_7_124_inst : DFFX1 port map( D => n1195, CLK => n4849, Q => 
                           RAM_7_124_port, QN => n_1928);
   RAM_reg_7_123_inst : DFFX1 port map( D => n1194, CLK => n4850, Q => 
                           RAM_7_123_port, QN => n_1929);
   RAM_reg_7_122_inst : DFFX1 port map( D => n1193, CLK => n4850, Q => 
                           RAM_7_122_port, QN => n_1930);
   RAM_reg_7_121_inst : DFFX1 port map( D => n1192, CLK => n4850, Q => 
                           RAM_7_121_port, QN => n_1931);
   RAM_reg_7_120_inst : DFFX1 port map( D => n1191, CLK => n4850, Q => 
                           RAM_7_120_port, QN => n_1932);
   RAM_reg_7_119_inst : DFFX1 port map( D => n1190, CLK => n4850, Q => 
                           RAM_7_119_port, QN => n_1933);
   RAM_reg_7_118_inst : DFFX1 port map( D => n1189, CLK => n4850, Q => 
                           RAM_7_118_port, QN => n_1934);
   RAM_reg_7_117_inst : DFFX1 port map( D => n1188, CLK => n4850, Q => 
                           RAM_7_117_port, QN => n_1935);
   RAM_reg_7_116_inst : DFFX1 port map( D => n1187, CLK => n4850, Q => 
                           RAM_7_116_port, QN => n_1936);
   RAM_reg_7_115_inst : DFFX1 port map( D => n1186, CLK => n4850, Q => 
                           RAM_7_115_port, QN => n_1937);
   RAM_reg_7_114_inst : DFFX1 port map( D => n1185, CLK => n4850, Q => 
                           RAM_7_114_port, QN => n_1938);
   RAM_reg_7_113_inst : DFFX1 port map( D => n1184, CLK => n4850, Q => 
                           RAM_7_113_port, QN => n_1939);
   RAM_reg_7_112_inst : DFFX1 port map( D => n1183, CLK => n4850, Q => 
                           RAM_7_112_port, QN => n_1940);
   RAM_reg_7_111_inst : DFFX1 port map( D => n1182, CLK => n4851, Q => 
                           RAM_7_111_port, QN => n_1941);
   RAM_reg_7_110_inst : DFFX1 port map( D => n1181, CLK => n4851, Q => 
                           RAM_7_110_port, QN => n_1942);
   RAM_reg_7_109_inst : DFFX1 port map( D => n1180, CLK => n4851, Q => 
                           RAM_7_109_port, QN => n_1943);
   RAM_reg_7_108_inst : DFFX1 port map( D => n1179, CLK => n4851, Q => 
                           RAM_7_108_port, QN => n_1944);
   RAM_reg_7_107_inst : DFFX1 port map( D => n1178, CLK => n4851, Q => 
                           RAM_7_107_port, QN => n_1945);
   RAM_reg_7_106_inst : DFFX1 port map( D => n1177, CLK => n4851, Q => 
                           RAM_7_106_port, QN => n_1946);
   RAM_reg_7_105_inst : DFFX1 port map( D => n1176, CLK => n4851, Q => 
                           RAM_7_105_port, QN => n_1947);
   RAM_reg_7_104_inst : DFFX1 port map( D => n1175, CLK => n4851, Q => 
                           RAM_7_104_port, QN => n_1948);
   RAM_reg_7_103_inst : DFFX1 port map( D => n1174, CLK => n4851, Q => 
                           RAM_7_103_port, QN => n_1949);
   RAM_reg_7_102_inst : DFFX1 port map( D => n1173, CLK => n4851, Q => 
                           RAM_7_102_port, QN => n_1950);
   RAM_reg_7_101_inst : DFFX1 port map( D => n1172, CLK => n4851, Q => 
                           RAM_7_101_port, QN => n_1951);
   RAM_reg_7_100_inst : DFFX1 port map( D => n1171, CLK => n4851, Q => 
                           RAM_7_100_port, QN => n_1952);
   RAM_reg_7_99_inst : DFFX1 port map( D => n1170, CLK => n4852, Q => 
                           RAM_7_99_port, QN => n_1953);
   RAM_reg_7_98_inst : DFFX1 port map( D => n1169, CLK => n4852, Q => 
                           RAM_7_98_port, QN => n_1954);
   RAM_reg_7_97_inst : DFFX1 port map( D => n1168, CLK => n4852, Q => 
                           RAM_7_97_port, QN => n_1955);
   RAM_reg_7_96_inst : DFFX1 port map( D => n1167, CLK => n4852, Q => 
                           RAM_7_96_port, QN => n_1956);
   RAM_reg_7_95_inst : DFFX1 port map( D => n1166, CLK => n4852, Q => 
                           RAM_7_95_port, QN => n_1957);
   RAM_reg_7_94_inst : DFFX1 port map( D => n1165, CLK => n4852, Q => 
                           RAM_7_94_port, QN => n_1958);
   RAM_reg_7_93_inst : DFFX1 port map( D => n1164, CLK => n4852, Q => 
                           RAM_7_93_port, QN => n_1959);
   RAM_reg_7_92_inst : DFFX1 port map( D => n1163, CLK => n4852, Q => 
                           RAM_7_92_port, QN => n_1960);
   RAM_reg_7_91_inst : DFFX1 port map( D => n1162, CLK => n4846, Q => 
                           RAM_7_91_port, QN => n_1961);
   RAM_reg_7_90_inst : DFFX1 port map( D => n1161, CLK => n4846, Q => 
                           RAM_7_90_port, QN => n_1962);
   RAM_reg_7_89_inst : DFFX1 port map( D => n1160, CLK => n4846, Q => 
                           RAM_7_89_port, QN => n_1963);
   RAM_reg_7_88_inst : DFFX1 port map( D => n1159, CLK => n4846, Q => 
                           RAM_7_88_port, QN => n_1964);
   RAM_reg_7_87_inst : DFFX1 port map( D => n1158, CLK => n4847, Q => 
                           RAM_7_87_port, QN => n_1965);
   RAM_reg_7_86_inst : DFFX1 port map( D => n1157, CLK => n4847, Q => 
                           RAM_7_86_port, QN => n_1966);
   RAM_reg_7_85_inst : DFFX1 port map( D => n1156, CLK => n4847, Q => 
                           RAM_7_85_port, QN => n_1967);
   RAM_reg_7_84_inst : DFFX1 port map( D => n1155, CLK => n4847, Q => 
                           RAM_7_84_port, QN => n_1968);
   RAM_reg_7_83_inst : DFFX1 port map( D => n1154, CLK => n4847, Q => 
                           RAM_7_83_port, QN => n_1969);
   RAM_reg_7_82_inst : DFFX1 port map( D => n1153, CLK => n4847, Q => 
                           RAM_7_82_port, QN => n_1970);
   RAM_reg_7_81_inst : DFFX1 port map( D => n1152, CLK => n4847, Q => 
                           RAM_7_81_port, QN => n_1971);
   RAM_reg_7_80_inst : DFFX1 port map( D => n1151, CLK => n4847, Q => 
                           RAM_7_80_port, QN => n_1972);
   RAM_reg_7_79_inst : DFFX1 port map( D => n1150, CLK => n4847, Q => 
                           RAM_7_79_port, QN => n_1973);
   RAM_reg_7_78_inst : DFFX1 port map( D => n1149, CLK => n4847, Q => 
                           RAM_7_78_port, QN => n_1974);
   RAM_reg_7_77_inst : DFFX1 port map( D => n1148, CLK => n4847, Q => 
                           RAM_7_77_port, QN => n_1975);
   RAM_reg_7_76_inst : DFFX1 port map( D => n1147, CLK => n4847, Q => 
                           RAM_7_76_port, QN => n_1976);
   RAM_reg_7_75_inst : DFFX1 port map( D => n1146, CLK => n4848, Q => 
                           RAM_7_75_port, QN => n_1977);
   RAM_reg_7_74_inst : DFFX1 port map( D => n1145, CLK => n4848, Q => 
                           RAM_7_74_port, QN => n_1978);
   RAM_reg_7_73_inst : DFFX1 port map( D => n1144, CLK => n4848, Q => 
                           RAM_7_73_port, QN => n_1979);
   RAM_reg_7_72_inst : DFFX1 port map( D => n1143, CLK => n4848, Q => 
                           RAM_7_72_port, QN => n_1980);
   RAM_reg_7_71_inst : DFFX1 port map( D => n1142, CLK => n4848, Q => 
                           RAM_7_71_port, QN => n_1981);
   RAM_reg_7_70_inst : DFFX1 port map( D => n1141, CLK => n4848, Q => 
                           RAM_7_70_port, QN => n_1982);
   RAM_reg_7_69_inst : DFFX1 port map( D => n1140, CLK => n4848, Q => 
                           RAM_7_69_port, QN => n_1983);
   RAM_reg_7_68_inst : DFFX1 port map( D => n1139, CLK => n4848, Q => 
                           RAM_7_68_port, QN => n_1984);
   RAM_reg_7_67_inst : DFFX1 port map( D => n1138, CLK => n4848, Q => 
                           RAM_7_67_port, QN => n_1985);
   RAM_reg_7_66_inst : DFFX1 port map( D => n1137, CLK => n4848, Q => 
                           RAM_7_66_port, QN => n_1986);
   RAM_reg_7_65_inst : DFFX1 port map( D => n1136, CLK => n4848, Q => 
                           RAM_7_65_port, QN => n_1987);
   RAM_reg_7_64_inst : DFFX1 port map( D => n1135, CLK => n4848, Q => 
                           RAM_7_64_port, QN => n_1988);
   RAM_reg_7_63_inst : DFFX1 port map( D => n1134, CLK => n4849, Q => 
                           RAM_7_63_port, QN => n_1989);
   RAM_reg_7_62_inst : DFFX1 port map( D => n1133, CLK => n4849, Q => 
                           RAM_7_62_port, QN => n_1990);
   RAM_reg_7_61_inst : DFFX1 port map( D => n1132, CLK => n4849, Q => 
                           RAM_7_61_port, QN => n_1991);
   RAM_reg_7_60_inst : DFFX1 port map( D => n1131, CLK => n4849, Q => 
                           RAM_7_60_port, QN => n_1992);
   RAM_reg_7_59_inst : DFFX1 port map( D => n1130, CLK => n4849, Q => 
                           RAM_7_59_port, QN => n_1993);
   RAM_reg_7_58_inst : DFFX1 port map( D => n1129, CLK => n4849, Q => 
                           RAM_7_58_port, QN => n_1994);
   RAM_reg_7_57_inst : DFFX1 port map( D => n1128, CLK => n4849, Q => 
                           RAM_7_57_port, QN => n_1995);
   RAM_reg_7_56_inst : DFFX1 port map( D => n1127, CLK => n4849, Q => 
                           RAM_7_56_port, QN => n_1996);
   RAM_reg_7_55_inst : DFFX1 port map( D => n1126, CLK => n4861, Q => 
                           RAM_7_55_port, QN => n_1997);
   RAM_reg_7_54_inst : DFFX1 port map( D => n1125, CLK => n4861, Q => 
                           RAM_7_54_port, QN => n_1998);
   RAM_reg_7_53_inst : DFFX1 port map( D => n1124, CLK => n4861, Q => 
                           RAM_7_53_port, QN => n_1999);
   RAM_reg_7_52_inst : DFFX1 port map( D => n1123, CLK => n4861, Q => 
                           RAM_7_52_port, QN => n_2000);
   RAM_reg_7_51_inst : DFFX1 port map( D => n1122, CLK => n4862, Q => 
                           RAM_7_51_port, QN => n_2001);
   RAM_reg_7_50_inst : DFFX1 port map( D => n1121, CLK => n4862, Q => 
                           RAM_7_50_port, QN => n_2002);
   RAM_reg_7_49_inst : DFFX1 port map( D => n1120, CLK => n4862, Q => 
                           RAM_7_49_port, QN => n_2003);
   RAM_reg_7_48_inst : DFFX1 port map( D => n1119, CLK => n4862, Q => 
                           RAM_7_48_port, QN => n_2004);
   RAM_reg_7_47_inst : DFFX1 port map( D => n1118, CLK => n4862, Q => 
                           RAM_7_47_port, QN => n_2005);
   RAM_reg_7_46_inst : DFFX1 port map( D => n1117, CLK => n4862, Q => 
                           RAM_7_46_port, QN => n_2006);
   RAM_reg_7_45_inst : DFFX1 port map( D => n1116, CLK => n4862, Q => 
                           RAM_7_45_port, QN => n_2007);
   RAM_reg_7_44_inst : DFFX1 port map( D => n1115, CLK => n4862, Q => 
                           RAM_7_44_port, QN => n_2008);
   RAM_reg_7_43_inst : DFFX1 port map( D => n1114, CLK => n4862, Q => 
                           RAM_7_43_port, QN => n_2009);
   RAM_reg_7_42_inst : DFFX1 port map( D => n1113, CLK => n4862, Q => 
                           RAM_7_42_port, QN => n_2010);
   RAM_reg_7_41_inst : DFFX1 port map( D => n1112, CLK => n4862, Q => 
                           RAM_7_41_port, QN => n_2011);
   RAM_reg_7_40_inst : DFFX1 port map( D => n1111, CLK => n4862, Q => 
                           RAM_7_40_port, QN => n_2012);
   RAM_reg_7_39_inst : DFFX1 port map( D => n1110, CLK => n4863, Q => 
                           RAM_7_39_port, QN => n_2013);
   RAM_reg_7_38_inst : DFFX1 port map( D => n1109, CLK => n4863, Q => 
                           RAM_7_38_port, QN => n_2014);
   RAM_reg_7_37_inst : DFFX1 port map( D => n1108, CLK => n4863, Q => 
                           RAM_7_37_port, QN => n_2015);
   RAM_reg_7_36_inst : DFFX1 port map( D => n1107, CLK => n4863, Q => 
                           RAM_7_36_port, QN => n_2016);
   RAM_reg_7_35_inst : DFFX1 port map( D => n1106, CLK => n4863, Q => 
                           RAM_7_35_port, QN => n_2017);
   RAM_reg_7_34_inst : DFFX1 port map( D => n1105, CLK => n4863, Q => 
                           RAM_7_34_port, QN => n_2018);
   RAM_reg_7_33_inst : DFFX1 port map( D => n1104, CLK => n4863, Q => 
                           RAM_7_33_port, QN => n_2019);
   RAM_reg_7_32_inst : DFFX1 port map( D => n1103, CLK => n4863, Q => 
                           RAM_7_32_port, QN => n_2020);
   RAM_reg_7_31_inst : DFFX1 port map( D => n1102, CLK => n4863, Q => 
                           RAM_7_31_port, QN => n_2021);
   RAM_reg_7_30_inst : DFFX1 port map( D => n1101, CLK => n4863, Q => 
                           RAM_7_30_port, QN => n_2022);
   RAM_reg_7_29_inst : DFFX1 port map( D => n1100, CLK => n4863, Q => 
                           RAM_7_29_port, QN => n_2023);
   RAM_reg_7_28_inst : DFFX1 port map( D => n1099, CLK => n4863, Q => 
                           RAM_7_28_port, QN => n_2024);
   RAM_reg_7_27_inst : DFFX1 port map( D => n1098, CLK => n4864, Q => 
                           RAM_7_27_port, QN => n_2025);
   RAM_reg_7_26_inst : DFFX1 port map( D => n1097, CLK => n4864, Q => 
                           RAM_7_26_port, QN => n_2026);
   RAM_reg_7_25_inst : DFFX1 port map( D => n1096, CLK => n4864, Q => 
                           RAM_7_25_port, QN => n_2027);
   RAM_reg_7_24_inst : DFFX1 port map( D => n1095, CLK => n4864, Q => 
                           RAM_7_24_port, QN => n_2028);
   RAM_reg_7_23_inst : DFFX1 port map( D => n1094, CLK => n4864, Q => 
                           RAM_7_23_port, QN => n_2029);
   RAM_reg_7_22_inst : DFFX1 port map( D => n1093, CLK => n4864, Q => 
                           RAM_7_22_port, QN => n_2030);
   RAM_reg_7_21_inst : DFFX1 port map( D => n1092, CLK => n4864, Q => 
                           RAM_7_21_port, QN => n_2031);
   RAM_reg_7_20_inst : DFFX1 port map( D => n1091, CLK => n4864, Q => 
                           RAM_7_20_port, QN => n_2032);
   RAM_reg_7_19_inst : DFFX1 port map( D => n1090, CLK => n4858, Q => 
                           RAM_7_19_port, QN => n_2033);
   RAM_reg_7_18_inst : DFFX1 port map( D => n1089, CLK => n4858, Q => 
                           RAM_7_18_port, QN => n_2034);
   RAM_reg_7_17_inst : DFFX1 port map( D => n1088, CLK => n4858, Q => 
                           RAM_7_17_port, QN => n_2035);
   RAM_reg_7_16_inst : DFFX1 port map( D => n1087, CLK => n4858, Q => 
                           RAM_7_16_port, QN => n_2036);
   RAM_reg_7_15_inst : DFFX1 port map( D => n1086, CLK => n4859, Q => 
                           RAM_7_15_port, QN => n_2037);
   RAM_reg_7_14_inst : DFFX1 port map( D => n1085, CLK => n4859, Q => 
                           RAM_7_14_port, QN => n_2038);
   RAM_reg_7_13_inst : DFFX1 port map( D => n1084, CLK => n4859, Q => 
                           RAM_7_13_port, QN => n_2039);
   RAM_reg_7_12_inst : DFFX1 port map( D => n1083, CLK => n4859, Q => 
                           RAM_7_12_port, QN => n_2040);
   RAM_reg_7_11_inst : DFFX1 port map( D => n1082, CLK => n4859, Q => 
                           RAM_7_11_port, QN => n_2041);
   RAM_reg_7_10_inst : DFFX1 port map( D => n1081, CLK => n4859, Q => 
                           RAM_7_10_port, QN => n_2042);
   RAM_reg_7_9_inst : DFFX1 port map( D => n1080, CLK => n4859, Q => 
                           RAM_7_9_port, QN => n_2043);
   RAM_reg_7_8_inst : DFFX1 port map( D => n1079, CLK => n4859, Q => 
                           RAM_7_8_port, QN => n_2044);
   RAM_reg_7_7_inst : DFFX1 port map( D => n1078, CLK => n4859, Q => 
                           RAM_7_7_port, QN => n_2045);
   RAM_reg_7_6_inst : DFFX1 port map( D => n1077, CLK => n4859, Q => 
                           RAM_7_6_port, QN => n_2046);
   RAM_reg_7_5_inst : DFFX1 port map( D => n1076, CLK => n4859, Q => 
                           RAM_7_5_port, QN => n_2047);
   RAM_reg_7_4_inst : DFFX1 port map( D => n1075, CLK => n4859, Q => 
                           RAM_7_4_port, QN => n_2048);
   RAM_reg_7_3_inst : DFFX1 port map( D => n1074, CLK => n4860, Q => 
                           RAM_7_3_port, QN => n_2049);
   RAM_reg_7_2_inst : DFFX1 port map( D => n1073, CLK => n4860, Q => 
                           RAM_7_2_port, QN => n_2050);
   RAM_reg_7_1_inst : DFFX1 port map( D => n1072, CLK => n4860, Q => 
                           RAM_7_1_port, QN => n_2051);
   RAM_reg_7_0_inst : DFFX1 port map( D => n1071, CLK => n4860, Q => 
                           RAM_7_0_port, QN => n_2052);
   RAM_reg_8_127_inst : DFFX1 port map( D => n1070, CLK => n4860, Q => 
                           RAM_8_127_port, QN => n_2053);
   RAM_reg_8_126_inst : DFFX1 port map( D => n1069, CLK => n4860, Q => 
                           RAM_8_126_port, QN => n_2054);
   RAM_reg_8_125_inst : DFFX1 port map( D => n1068, CLK => n4860, Q => 
                           RAM_8_125_port, QN => n_2055);
   RAM_reg_8_124_inst : DFFX1 port map( D => n1067, CLK => n4860, Q => 
                           RAM_8_124_port, QN => n_2056);
   RAM_reg_8_123_inst : DFFX1 port map( D => n1066, CLK => n4860, Q => 
                           RAM_8_123_port, QN => n_2057);
   RAM_reg_8_122_inst : DFFX1 port map( D => n1065, CLK => n4860, Q => 
                           RAM_8_122_port, QN => n_2058);
   RAM_reg_8_121_inst : DFFX1 port map( D => n1064, CLK => n4860, Q => 
                           RAM_8_121_port, QN => n_2059);
   RAM_reg_8_120_inst : DFFX1 port map( D => n1063, CLK => n4860, Q => 
                           RAM_8_120_port, QN => n_2060);
   RAM_reg_8_119_inst : DFFX1 port map( D => n1062, CLK => n4861, Q => 
                           RAM_8_119_port, QN => n_2061);
   RAM_reg_8_118_inst : DFFX1 port map( D => n1061, CLK => n4861, Q => 
                           RAM_8_118_port, QN => n_2062);
   RAM_reg_8_117_inst : DFFX1 port map( D => n1060, CLK => n4861, Q => 
                           RAM_8_117_port, QN => n_2063);
   RAM_reg_8_116_inst : DFFX1 port map( D => n1059, CLK => n4861, Q => 
                           RAM_8_116_port, QN => n_2064);
   RAM_reg_8_115_inst : DFFX1 port map( D => n1058, CLK => n4861, Q => 
                           RAM_8_115_port, QN => n_2065);
   RAM_reg_8_114_inst : DFFX1 port map( D => n1057, CLK => n4861, Q => 
                           RAM_8_114_port, QN => n_2066);
   RAM_reg_8_113_inst : DFFX1 port map( D => n1056, CLK => n4861, Q => 
                           RAM_8_113_port, QN => n_2067);
   RAM_reg_8_112_inst : DFFX1 port map( D => n1055, CLK => n4861, Q => 
                           RAM_8_112_port, QN => n_2068);
   RAM_reg_8_111_inst : DFFX1 port map( D => n1054, CLK => n4855, Q => 
                           RAM_8_111_port, QN => n_2069);
   RAM_reg_8_110_inst : DFFX1 port map( D => n1053, CLK => n4855, Q => 
                           RAM_8_110_port, QN => n_2070);
   RAM_reg_8_109_inst : DFFX1 port map( D => n1052, CLK => n4855, Q => 
                           RAM_8_109_port, QN => n_2071);
   RAM_reg_8_108_inst : DFFX1 port map( D => n1051, CLK => n4855, Q => 
                           RAM_8_108_port, QN => n_2072);
   RAM_reg_8_107_inst : DFFX1 port map( D => n1050, CLK => n4856, Q => 
                           RAM_8_107_port, QN => n_2073);
   RAM_reg_8_106_inst : DFFX1 port map( D => n1049, CLK => n4856, Q => 
                           RAM_8_106_port, QN => n_2074);
   RAM_reg_8_105_inst : DFFX1 port map( D => n1048, CLK => n4856, Q => 
                           RAM_8_105_port, QN => n_2075);
   RAM_reg_8_104_inst : DFFX1 port map( D => n1047, CLK => n4856, Q => 
                           RAM_8_104_port, QN => n_2076);
   RAM_reg_8_103_inst : DFFX1 port map( D => n1046, CLK => n4856, Q => 
                           RAM_8_103_port, QN => n_2077);
   RAM_reg_8_102_inst : DFFX1 port map( D => n1045, CLK => n4856, Q => 
                           RAM_8_102_port, QN => n_2078);
   RAM_reg_8_101_inst : DFFX1 port map( D => n1044, CLK => n4856, Q => 
                           RAM_8_101_port, QN => n_2079);
   RAM_reg_8_100_inst : DFFX1 port map( D => n1043, CLK => n4856, Q => 
                           RAM_8_100_port, QN => n_2080);
   RAM_reg_8_99_inst : DFFX1 port map( D => n1042, CLK => n4856, Q => 
                           RAM_8_99_port, QN => n_2081);
   RAM_reg_8_98_inst : DFFX1 port map( D => n1041, CLK => n4856, Q => 
                           RAM_8_98_port, QN => n_2082);
   RAM_reg_8_97_inst : DFFX1 port map( D => n1040, CLK => n4856, Q => 
                           RAM_8_97_port, QN => n_2083);
   RAM_reg_8_96_inst : DFFX1 port map( D => n1039, CLK => n4856, Q => 
                           RAM_8_96_port, QN => n_2084);
   RAM_reg_8_95_inst : DFFX1 port map( D => n1038, CLK => n4857, Q => 
                           RAM_8_95_port, QN => n_2085);
   RAM_reg_8_94_inst : DFFX1 port map( D => n1037, CLK => n4857, Q => 
                           RAM_8_94_port, QN => n_2086);
   RAM_reg_8_93_inst : DFFX1 port map( D => n1036, CLK => n4857, Q => 
                           RAM_8_93_port, QN => n_2087);
   RAM_reg_8_92_inst : DFFX1 port map( D => n1035, CLK => n4857, Q => 
                           RAM_8_92_port, QN => n_2088);
   RAM_reg_8_91_inst : DFFX1 port map( D => n1034, CLK => n4857, Q => 
                           RAM_8_91_port, QN => n_2089);
   RAM_reg_8_90_inst : DFFX1 port map( D => n1033, CLK => n4857, Q => 
                           RAM_8_90_port, QN => n_2090);
   RAM_reg_8_89_inst : DFFX1 port map( D => n1032, CLK => n4857, Q => 
                           RAM_8_89_port, QN => n_2091);
   RAM_reg_8_88_inst : DFFX1 port map( D => n1031, CLK => n4857, Q => 
                           RAM_8_88_port, QN => n_2092);
   RAM_reg_8_87_inst : DFFX1 port map( D => n1030, CLK => n4857, Q => 
                           RAM_8_87_port, QN => n_2093);
   RAM_reg_8_86_inst : DFFX1 port map( D => n1029, CLK => n4857, Q => 
                           RAM_8_86_port, QN => n_2094);
   RAM_reg_8_85_inst : DFFX1 port map( D => n1028, CLK => n4857, Q => 
                           RAM_8_85_port, QN => n_2095);
   RAM_reg_8_84_inst : DFFX1 port map( D => n1027, CLK => n4857, Q => 
                           RAM_8_84_port, QN => n_2096);
   RAM_reg_8_83_inst : DFFX1 port map( D => n1026, CLK => n4858, Q => 
                           RAM_8_83_port, QN => n_2097);
   RAM_reg_8_82_inst : DFFX1 port map( D => n1025, CLK => n4858, Q => 
                           RAM_8_82_port, QN => n_2098);
   RAM_reg_8_81_inst : DFFX1 port map( D => n1024, CLK => n4858, Q => 
                           RAM_8_81_port, QN => n_2099);
   RAM_reg_8_80_inst : DFFX1 port map( D => n1023, CLK => n4858, Q => 
                           RAM_8_80_port, QN => n_2100);
   RAM_reg_8_79_inst : DFFX1 port map( D => n1022, CLK => n4858, Q => 
                           RAM_8_79_port, QN => n_2101);
   RAM_reg_8_78_inst : DFFX1 port map( D => n1021, CLK => n4858, Q => 
                           RAM_8_78_port, QN => n_2102);
   RAM_reg_8_77_inst : DFFX1 port map( D => n1020, CLK => n4858, Q => 
                           RAM_8_77_port, QN => n_2103);
   RAM_reg_8_76_inst : DFFX1 port map( D => n1019, CLK => n4858, Q => 
                           RAM_8_76_port, QN => n_2104);
   RAM_reg_8_75_inst : DFFX1 port map( D => n1018, CLK => n4870, Q => 
                           RAM_8_75_port, QN => n_2105);
   RAM_reg_8_74_inst : DFFX1 port map( D => n1017, CLK => n4870, Q => 
                           RAM_8_74_port, QN => n_2106);
   RAM_reg_8_73_inst : DFFX1 port map( D => n1016, CLK => n4870, Q => 
                           RAM_8_73_port, QN => n_2107);
   RAM_reg_8_72_inst : DFFX1 port map( D => n1015, CLK => n4870, Q => 
                           RAM_8_72_port, QN => n_2108);
   RAM_reg_8_71_inst : DFFX1 port map( D => n1014, CLK => n4871, Q => 
                           RAM_8_71_port, QN => n_2109);
   RAM_reg_8_70_inst : DFFX1 port map( D => n1013, CLK => n4871, Q => 
                           RAM_8_70_port, QN => n_2110);
   RAM_reg_8_69_inst : DFFX1 port map( D => n1012, CLK => n4871, Q => 
                           RAM_8_69_port, QN => n_2111);
   RAM_reg_8_68_inst : DFFX1 port map( D => n1011, CLK => n4871, Q => 
                           RAM_8_68_port, QN => n_2112);
   RAM_reg_8_67_inst : DFFX1 port map( D => n1010, CLK => n4871, Q => 
                           RAM_8_67_port, QN => n_2113);
   RAM_reg_8_66_inst : DFFX1 port map( D => n1009, CLK => n4871, Q => 
                           RAM_8_66_port, QN => n_2114);
   RAM_reg_8_65_inst : DFFX1 port map( D => n1008, CLK => n4871, Q => 
                           RAM_8_65_port, QN => n_2115);
   RAM_reg_8_64_inst : DFFX1 port map( D => n1007, CLK => n4871, Q => 
                           RAM_8_64_port, QN => n_2116);
   RAM_reg_8_63_inst : DFFX1 port map( D => n1006, CLK => n4871, Q => 
                           RAM_8_63_port, QN => n_2117);
   RAM_reg_8_62_inst : DFFX1 port map( D => n1005, CLK => n4871, Q => 
                           RAM_8_62_port, QN => n_2118);
   RAM_reg_8_61_inst : DFFX1 port map( D => n1004, CLK => n4871, Q => 
                           RAM_8_61_port, QN => n_2119);
   RAM_reg_8_60_inst : DFFX1 port map( D => n1003, CLK => n4871, Q => 
                           RAM_8_60_port, QN => n_2120);
   RAM_reg_8_59_inst : DFFX1 port map( D => n1002, CLK => n4872, Q => 
                           RAM_8_59_port, QN => n_2121);
   RAM_reg_8_58_inst : DFFX1 port map( D => n1001, CLK => n4872, Q => 
                           RAM_8_58_port, QN => n_2122);
   RAM_reg_8_57_inst : DFFX1 port map( D => n1000, CLK => n4872, Q => 
                           RAM_8_57_port, QN => n_2123);
   RAM_reg_8_56_inst : DFFX1 port map( D => n999, CLK => n4872, Q => 
                           RAM_8_56_port, QN => n_2124);
   RAM_reg_8_55_inst : DFFX1 port map( D => n998, CLK => n4872, Q => 
                           RAM_8_55_port, QN => n_2125);
   RAM_reg_8_54_inst : DFFX1 port map( D => n997, CLK => n4872, Q => 
                           RAM_8_54_port, QN => n_2126);
   RAM_reg_8_53_inst : DFFX1 port map( D => n996, CLK => n4872, Q => 
                           RAM_8_53_port, QN => n_2127);
   RAM_reg_8_52_inst : DFFX1 port map( D => n995, CLK => n4872, Q => 
                           RAM_8_52_port, QN => n_2128);
   RAM_reg_8_51_inst : DFFX1 port map( D => n994, CLK => n4872, Q => 
                           RAM_8_51_port, QN => n_2129);
   RAM_reg_8_50_inst : DFFX1 port map( D => n993, CLK => n4872, Q => 
                           RAM_8_50_port, QN => n_2130);
   RAM_reg_8_49_inst : DFFX1 port map( D => n992, CLK => n4872, Q => 
                           RAM_8_49_port, QN => n_2131);
   RAM_reg_8_48_inst : DFFX1 port map( D => n991, CLK => n4872, Q => 
                           RAM_8_48_port, QN => n_2132);
   RAM_reg_8_47_inst : DFFX1 port map( D => n990, CLK => n4873, Q => 
                           RAM_8_47_port, QN => n_2133);
   RAM_reg_8_46_inst : DFFX1 port map( D => n989, CLK => n4873, Q => 
                           RAM_8_46_port, QN => n_2134);
   RAM_reg_8_45_inst : DFFX1 port map( D => n988, CLK => n4873, Q => 
                           RAM_8_45_port, QN => n_2135);
   RAM_reg_8_44_inst : DFFX1 port map( D => n987, CLK => n4873, Q => 
                           RAM_8_44_port, QN => n_2136);
   RAM_reg_8_43_inst : DFFX1 port map( D => n986, CLK => n4873, Q => 
                           RAM_8_43_port, QN => n_2137);
   RAM_reg_8_42_inst : DFFX1 port map( D => n985, CLK => n4873, Q => 
                           RAM_8_42_port, QN => n_2138);
   RAM_reg_8_41_inst : DFFX1 port map( D => n984, CLK => n4873, Q => 
                           RAM_8_41_port, QN => n_2139);
   RAM_reg_8_40_inst : DFFX1 port map( D => n983, CLK => n4873, Q => 
                           RAM_8_40_port, QN => n_2140);
   RAM_reg_8_39_inst : DFFX1 port map( D => n982, CLK => n4867, Q => 
                           RAM_8_39_port, QN => n_2141);
   RAM_reg_8_38_inst : DFFX1 port map( D => n981, CLK => n4867, Q => 
                           RAM_8_38_port, QN => n_2142);
   RAM_reg_8_37_inst : DFFX1 port map( D => n980, CLK => n4867, Q => 
                           RAM_8_37_port, QN => n_2143);
   RAM_reg_8_36_inst : DFFX1 port map( D => n979, CLK => n4867, Q => 
                           RAM_8_36_port, QN => n_2144);
   RAM_reg_8_35_inst : DFFX1 port map( D => n978, CLK => n4868, Q => 
                           RAM_8_35_port, QN => n_2145);
   RAM_reg_8_34_inst : DFFX1 port map( D => n977, CLK => n4868, Q => 
                           RAM_8_34_port, QN => n_2146);
   RAM_reg_8_33_inst : DFFX1 port map( D => n976, CLK => n4868, Q => 
                           RAM_8_33_port, QN => n_2147);
   RAM_reg_8_32_inst : DFFX1 port map( D => n975, CLK => n4868, Q => 
                           RAM_8_32_port, QN => n_2148);
   RAM_reg_8_31_inst : DFFX1 port map( D => n974, CLK => n4868, Q => 
                           RAM_8_31_port, QN => n_2149);
   RAM_reg_8_30_inst : DFFX1 port map( D => n973, CLK => n4868, Q => 
                           RAM_8_30_port, QN => n_2150);
   RAM_reg_8_29_inst : DFFX1 port map( D => n972, CLK => n4868, Q => 
                           RAM_8_29_port, QN => n_2151);
   RAM_reg_8_28_inst : DFFX1 port map( D => n971, CLK => n4868, Q => 
                           RAM_8_28_port, QN => n_2152);
   RAM_reg_8_27_inst : DFFX1 port map( D => n970, CLK => n4868, Q => 
                           RAM_8_27_port, QN => n_2153);
   RAM_reg_8_26_inst : DFFX1 port map( D => n969, CLK => n4868, Q => 
                           RAM_8_26_port, QN => n_2154);
   RAM_reg_8_25_inst : DFFX1 port map( D => n968, CLK => n4868, Q => 
                           RAM_8_25_port, QN => n_2155);
   RAM_reg_8_24_inst : DFFX1 port map( D => n967, CLK => n4868, Q => 
                           RAM_8_24_port, QN => n_2156);
   RAM_reg_8_23_inst : DFFX1 port map( D => n966, CLK => n4869, Q => 
                           RAM_8_23_port, QN => n_2157);
   RAM_reg_8_22_inst : DFFX1 port map( D => n965, CLK => n4869, Q => 
                           RAM_8_22_port, QN => n_2158);
   RAM_reg_8_21_inst : DFFX1 port map( D => n964, CLK => n4869, Q => 
                           RAM_8_21_port, QN => n_2159);
   RAM_reg_8_20_inst : DFFX1 port map( D => n963, CLK => n4869, Q => 
                           RAM_8_20_port, QN => n_2160);
   RAM_reg_8_19_inst : DFFX1 port map( D => n962, CLK => n4869, Q => 
                           RAM_8_19_port, QN => n_2161);
   RAM_reg_8_18_inst : DFFX1 port map( D => n961, CLK => n4869, Q => 
                           RAM_8_18_port, QN => n_2162);
   RAM_reg_8_17_inst : DFFX1 port map( D => n960, CLK => n4869, Q => 
                           RAM_8_17_port, QN => n_2163);
   RAM_reg_8_16_inst : DFFX1 port map( D => n959, CLK => n4869, Q => 
                           RAM_8_16_port, QN => n_2164);
   RAM_reg_8_15_inst : DFFX1 port map( D => n958, CLK => n4869, Q => 
                           RAM_8_15_port, QN => n_2165);
   RAM_reg_8_14_inst : DFFX1 port map( D => n957, CLK => n4869, Q => 
                           RAM_8_14_port, QN => n_2166);
   RAM_reg_8_13_inst : DFFX1 port map( D => n956, CLK => n4869, Q => 
                           RAM_8_13_port, QN => n_2167);
   RAM_reg_8_12_inst : DFFX1 port map( D => n955, CLK => n4869, Q => 
                           RAM_8_12_port, QN => n_2168);
   RAM_reg_8_11_inst : DFFX1 port map( D => n954, CLK => n4870, Q => 
                           RAM_8_11_port, QN => n_2169);
   RAM_reg_8_10_inst : DFFX1 port map( D => n953, CLK => n4870, Q => 
                           RAM_8_10_port, QN => n_2170);
   RAM_reg_8_9_inst : DFFX1 port map( D => n952, CLK => n4870, Q => 
                           RAM_8_9_port, QN => n_2171);
   RAM_reg_8_8_inst : DFFX1 port map( D => n951, CLK => n4870, Q => 
                           RAM_8_8_port, QN => n_2172);
   RAM_reg_8_7_inst : DFFX1 port map( D => n950, CLK => n4870, Q => 
                           RAM_8_7_port, QN => n_2173);
   RAM_reg_8_6_inst : DFFX1 port map( D => n949, CLK => n4870, Q => 
                           RAM_8_6_port, QN => n_2174);
   RAM_reg_8_5_inst : DFFX1 port map( D => n948, CLK => n4870, Q => 
                           RAM_8_5_port, QN => n_2175);
   RAM_reg_8_4_inst : DFFX1 port map( D => n947, CLK => n4870, Q => 
                           RAM_8_4_port, QN => n_2176);
   RAM_reg_8_3_inst : DFFX1 port map( D => n946, CLK => n4864, Q => 
                           RAM_8_3_port, QN => n_2177);
   RAM_reg_8_2_inst : DFFX1 port map( D => n945, CLK => n4864, Q => 
                           RAM_8_2_port, QN => n_2178);
   RAM_reg_8_1_inst : DFFX1 port map( D => n944, CLK => n4864, Q => 
                           RAM_8_1_port, QN => n_2179);
   RAM_reg_8_0_inst : DFFX1 port map( D => n943, CLK => n4864, Q => 
                           RAM_8_0_port, QN => n_2180);
   RAM_reg_9_127_inst : DFFX1 port map( D => n942, CLK => n4865, Q => 
                           RAM_9_127_port, QN => n_2181);
   RAM_reg_9_126_inst : DFFX1 port map( D => n941, CLK => n4865, Q => 
                           RAM_9_126_port, QN => n_2182);
   RAM_reg_9_125_inst : DFFX1 port map( D => n940, CLK => n4865, Q => 
                           RAM_9_125_port, QN => n_2183);
   RAM_reg_9_124_inst : DFFX1 port map( D => n939, CLK => n4865, Q => 
                           RAM_9_124_port, QN => n_2184);
   RAM_reg_9_123_inst : DFFX1 port map( D => n938, CLK => n4865, Q => 
                           RAM_9_123_port, QN => n_2185);
   RAM_reg_9_122_inst : DFFX1 port map( D => n937, CLK => n4865, Q => 
                           RAM_9_122_port, QN => n_2186);
   RAM_reg_9_121_inst : DFFX1 port map( D => n936, CLK => n4865, Q => 
                           RAM_9_121_port, QN => n_2187);
   RAM_reg_9_120_inst : DFFX1 port map( D => n935, CLK => n4865, Q => 
                           RAM_9_120_port, QN => n_2188);
   RAM_reg_9_119_inst : DFFX1 port map( D => n934, CLK => n4865, Q => 
                           RAM_9_119_port, QN => n_2189);
   RAM_reg_9_118_inst : DFFX1 port map( D => n933, CLK => n4865, Q => 
                           RAM_9_118_port, QN => n_2190);
   RAM_reg_9_117_inst : DFFX1 port map( D => n932, CLK => n4865, Q => 
                           RAM_9_117_port, QN => n_2191);
   RAM_reg_9_116_inst : DFFX1 port map( D => n931, CLK => n4865, Q => 
                           RAM_9_116_port, QN => n_2192);
   RAM_reg_9_115_inst : DFFX1 port map( D => n930, CLK => n4866, Q => 
                           RAM_9_115_port, QN => n_2193);
   RAM_reg_9_114_inst : DFFX1 port map( D => n929, CLK => n4866, Q => 
                           RAM_9_114_port, QN => n_2194);
   RAM_reg_9_113_inst : DFFX1 port map( D => n928, CLK => n4866, Q => 
                           RAM_9_113_port, QN => n_2195);
   RAM_reg_9_112_inst : DFFX1 port map( D => n927, CLK => n4866, Q => 
                           RAM_9_112_port, QN => n_2196);
   RAM_reg_9_111_inst : DFFX1 port map( D => n926, CLK => n4866, Q => 
                           RAM_9_111_port, QN => n_2197);
   RAM_reg_9_110_inst : DFFX1 port map( D => n925, CLK => n4866, Q => 
                           RAM_9_110_port, QN => n_2198);
   RAM_reg_9_109_inst : DFFX1 port map( D => n924, CLK => n4866, Q => 
                           RAM_9_109_port, QN => n_2199);
   RAM_reg_9_108_inst : DFFX1 port map( D => n923, CLK => n4866, Q => 
                           RAM_9_108_port, QN => n_2200);
   RAM_reg_9_107_inst : DFFX1 port map( D => n922, CLK => n4866, Q => 
                           RAM_9_107_port, QN => n_2201);
   RAM_reg_9_106_inst : DFFX1 port map( D => n921, CLK => n4866, Q => 
                           RAM_9_106_port, QN => n_2202);
   RAM_reg_9_105_inst : DFFX1 port map( D => n920, CLK => n4866, Q => 
                           RAM_9_105_port, QN => n_2203);
   RAM_reg_9_104_inst : DFFX1 port map( D => n919, CLK => n4866, Q => 
                           RAM_9_104_port, QN => n_2204);
   RAM_reg_9_103_inst : DFFX1 port map( D => n918, CLK => n4867, Q => 
                           RAM_9_103_port, QN => n_2205);
   RAM_reg_9_102_inst : DFFX1 port map( D => n917, CLK => n4867, Q => 
                           RAM_9_102_port, QN => n_2206);
   RAM_reg_9_101_inst : DFFX1 port map( D => n916, CLK => n4867, Q => 
                           RAM_9_101_port, QN => n_2207);
   RAM_reg_9_100_inst : DFFX1 port map( D => n915, CLK => n4867, Q => 
                           RAM_9_100_port, QN => n_2208);
   RAM_reg_9_99_inst : DFFX1 port map( D => n914, CLK => n4867, Q => 
                           RAM_9_99_port, QN => n_2209);
   RAM_reg_9_98_inst : DFFX1 port map( D => n913, CLK => n4867, Q => 
                           RAM_9_98_port, QN => n_2210);
   RAM_reg_9_97_inst : DFFX1 port map( D => n912, CLK => n4867, Q => 
                           RAM_9_97_port, QN => n_2211);
   RAM_reg_9_96_inst : DFFX1 port map( D => n911, CLK => n4867, Q => 
                           RAM_9_96_port, QN => n_2212);
   RAM_reg_9_95_inst : DFFX1 port map( D => n910, CLK => n4879, Q => 
                           RAM_9_95_port, QN => n_2213);
   RAM_reg_9_94_inst : DFFX1 port map( D => n909, CLK => n4879, Q => 
                           RAM_9_94_port, QN => n_2214);
   RAM_reg_9_93_inst : DFFX1 port map( D => n908, CLK => n4879, Q => 
                           RAM_9_93_port, QN => n_2215);
   RAM_reg_9_92_inst : DFFX1 port map( D => n907, CLK => n4879, Q => 
                           RAM_9_92_port, QN => n_2216);
   RAM_reg_9_91_inst : DFFX1 port map( D => n906, CLK => n4880, Q => 
                           RAM_9_91_port, QN => n_2217);
   RAM_reg_9_90_inst : DFFX1 port map( D => n905, CLK => n4880, Q => 
                           RAM_9_90_port, QN => n_2218);
   RAM_reg_9_89_inst : DFFX1 port map( D => n904, CLK => n4880, Q => 
                           RAM_9_89_port, QN => n_2219);
   RAM_reg_9_88_inst : DFFX1 port map( D => n903, CLK => n4880, Q => 
                           RAM_9_88_port, QN => n_2220);
   RAM_reg_9_87_inst : DFFX1 port map( D => n902, CLK => n4880, Q => 
                           RAM_9_87_port, QN => n_2221);
   RAM_reg_9_86_inst : DFFX1 port map( D => n901, CLK => n4880, Q => 
                           RAM_9_86_port, QN => n_2222);
   RAM_reg_9_85_inst : DFFX1 port map( D => n900, CLK => n4880, Q => 
                           RAM_9_85_port, QN => n_2223);
   RAM_reg_9_84_inst : DFFX1 port map( D => n899, CLK => n4880, Q => 
                           RAM_9_84_port, QN => n_2224);
   RAM_reg_9_83_inst : DFFX1 port map( D => n898, CLK => n4880, Q => 
                           RAM_9_83_port, QN => n_2225);
   RAM_reg_9_82_inst : DFFX1 port map( D => n897, CLK => n4880, Q => 
                           RAM_9_82_port, QN => n_2226);
   RAM_reg_9_81_inst : DFFX1 port map( D => n896, CLK => n4880, Q => 
                           RAM_9_81_port, QN => n_2227);
   RAM_reg_9_80_inst : DFFX1 port map( D => n895, CLK => n4880, Q => 
                           RAM_9_80_port, QN => n_2228);
   RAM_reg_9_79_inst : DFFX1 port map( D => n894, CLK => n4881, Q => 
                           RAM_9_79_port, QN => n_2229);
   RAM_reg_9_78_inst : DFFX1 port map( D => n893, CLK => n4881, Q => 
                           RAM_9_78_port, QN => n_2230);
   RAM_reg_9_77_inst : DFFX1 port map( D => n892, CLK => n4881, Q => 
                           RAM_9_77_port, QN => n_2231);
   RAM_reg_9_76_inst : DFFX1 port map( D => n891, CLK => n4881, Q => 
                           RAM_9_76_port, QN => n_2232);
   RAM_reg_9_75_inst : DFFX1 port map( D => n890, CLK => n4881, Q => 
                           RAM_9_75_port, QN => n_2233);
   RAM_reg_9_74_inst : DFFX1 port map( D => n889, CLK => n4881, Q => 
                           RAM_9_74_port, QN => n_2234);
   RAM_reg_9_73_inst : DFFX1 port map( D => n888, CLK => n4881, Q => 
                           RAM_9_73_port, QN => n_2235);
   RAM_reg_9_72_inst : DFFX1 port map( D => n887, CLK => n4881, Q => 
                           RAM_9_72_port, QN => n_2236);
   RAM_reg_9_71_inst : DFFX1 port map( D => n886, CLK => n4881, Q => 
                           RAM_9_71_port, QN => n_2237);
   RAM_reg_9_70_inst : DFFX1 port map( D => n885, CLK => n4881, Q => 
                           RAM_9_70_port, QN => n_2238);
   RAM_reg_9_69_inst : DFFX1 port map( D => n884, CLK => n4881, Q => 
                           RAM_9_69_port, QN => n_2239);
   RAM_reg_9_68_inst : DFFX1 port map( D => n883, CLK => n4881, Q => 
                           RAM_9_68_port, QN => n_2240);
   RAM_reg_9_67_inst : DFFX1 port map( D => n882, CLK => n4882, Q => 
                           RAM_9_67_port, QN => n_2241);
   RAM_reg_9_66_inst : DFFX1 port map( D => n881, CLK => n4882, Q => 
                           RAM_9_66_port, QN => n_2242);
   RAM_reg_9_65_inst : DFFX1 port map( D => n880, CLK => n4882, Q => 
                           RAM_9_65_port, QN => n_2243);
   RAM_reg_9_64_inst : DFFX1 port map( D => n879, CLK => n4882, Q => 
                           RAM_9_64_port, QN => n_2244);
   RAM_reg_9_63_inst : DFFX1 port map( D => n878, CLK => n4882, Q => 
                           RAM_9_63_port, QN => n_2245);
   RAM_reg_9_62_inst : DFFX1 port map( D => n877, CLK => n4882, Q => 
                           RAM_9_62_port, QN => n_2246);
   RAM_reg_9_61_inst : DFFX1 port map( D => n876, CLK => n4882, Q => 
                           RAM_9_61_port, QN => n_2247);
   RAM_reg_9_60_inst : DFFX1 port map( D => n875, CLK => n4882, Q => 
                           RAM_9_60_port, QN => n_2248);
   RAM_reg_9_59_inst : DFFX1 port map( D => n874, CLK => n4876, Q => 
                           RAM_9_59_port, QN => n_2249);
   RAM_reg_9_58_inst : DFFX1 port map( D => n873, CLK => n4876, Q => 
                           RAM_9_58_port, QN => n_2250);
   RAM_reg_9_57_inst : DFFX1 port map( D => n872, CLK => n4876, Q => 
                           RAM_9_57_port, QN => n_2251);
   RAM_reg_9_56_inst : DFFX1 port map( D => n871, CLK => n4876, Q => 
                           RAM_9_56_port, QN => n_2252);
   RAM_reg_9_55_inst : DFFX1 port map( D => n870, CLK => n4877, Q => 
                           RAM_9_55_port, QN => n_2253);
   RAM_reg_9_54_inst : DFFX1 port map( D => n869, CLK => n4877, Q => 
                           RAM_9_54_port, QN => n_2254);
   RAM_reg_9_53_inst : DFFX1 port map( D => n868, CLK => n4877, Q => 
                           RAM_9_53_port, QN => n_2255);
   RAM_reg_9_52_inst : DFFX1 port map( D => n867, CLK => n4877, Q => 
                           RAM_9_52_port, QN => n_2256);
   RAM_reg_9_51_inst : DFFX1 port map( D => n866, CLK => n4877, Q => 
                           RAM_9_51_port, QN => n_2257);
   RAM_reg_9_50_inst : DFFX1 port map( D => n865, CLK => n4877, Q => 
                           RAM_9_50_port, QN => n_2258);
   RAM_reg_9_49_inst : DFFX1 port map( D => n864, CLK => n4877, Q => 
                           RAM_9_49_port, QN => n_2259);
   RAM_reg_9_48_inst : DFFX1 port map( D => n863, CLK => n4877, Q => 
                           RAM_9_48_port, QN => n_2260);
   RAM_reg_9_47_inst : DFFX1 port map( D => n862, CLK => n4877, Q => 
                           RAM_9_47_port, QN => n_2261);
   RAM_reg_9_46_inst : DFFX1 port map( D => n861, CLK => n4877, Q => 
                           RAM_9_46_port, QN => n_2262);
   RAM_reg_9_45_inst : DFFX1 port map( D => n860, CLK => n4877, Q => 
                           RAM_9_45_port, QN => n_2263);
   RAM_reg_9_44_inst : DFFX1 port map( D => n859, CLK => n4877, Q => 
                           RAM_9_44_port, QN => n_2264);
   RAM_reg_9_43_inst : DFFX1 port map( D => n858, CLK => n4878, Q => 
                           RAM_9_43_port, QN => n_2265);
   RAM_reg_9_42_inst : DFFX1 port map( D => n857, CLK => n4878, Q => 
                           RAM_9_42_port, QN => n_2266);
   RAM_reg_9_41_inst : DFFX1 port map( D => n856, CLK => n4878, Q => 
                           RAM_9_41_port, QN => n_2267);
   RAM_reg_9_40_inst : DFFX1 port map( D => n855, CLK => n4878, Q => 
                           RAM_9_40_port, QN => n_2268);
   RAM_reg_9_39_inst : DFFX1 port map( D => n854, CLK => n4878, Q => 
                           RAM_9_39_port, QN => n_2269);
   RAM_reg_9_38_inst : DFFX1 port map( D => n853, CLK => n4878, Q => 
                           RAM_9_38_port, QN => n_2270);
   RAM_reg_9_37_inst : DFFX1 port map( D => n852, CLK => n4878, Q => 
                           RAM_9_37_port, QN => n_2271);
   RAM_reg_9_36_inst : DFFX1 port map( D => n851, CLK => n4878, Q => 
                           RAM_9_36_port, QN => n_2272);
   RAM_reg_9_35_inst : DFFX1 port map( D => n850, CLK => n4878, Q => 
                           RAM_9_35_port, QN => n_2273);
   RAM_reg_9_34_inst : DFFX1 port map( D => n849, CLK => n4878, Q => 
                           RAM_9_34_port, QN => n_2274);
   RAM_reg_9_33_inst : DFFX1 port map( D => n848, CLK => n4878, Q => 
                           RAM_9_33_port, QN => n_2275);
   RAM_reg_9_32_inst : DFFX1 port map( D => n847, CLK => n4878, Q => 
                           RAM_9_32_port, QN => n_2276);
   RAM_reg_9_31_inst : DFFX1 port map( D => n846, CLK => n4879, Q => 
                           RAM_9_31_port, QN => n_2277);
   RAM_reg_9_30_inst : DFFX1 port map( D => n845, CLK => n4879, Q => 
                           RAM_9_30_port, QN => n_2278);
   RAM_reg_9_29_inst : DFFX1 port map( D => n844, CLK => n4879, Q => 
                           RAM_9_29_port, QN => n_2279);
   RAM_reg_9_28_inst : DFFX1 port map( D => n843, CLK => n4879, Q => 
                           RAM_9_28_port, QN => n_2280);
   RAM_reg_9_27_inst : DFFX1 port map( D => n842, CLK => n4879, Q => 
                           RAM_9_27_port, QN => n_2281);
   RAM_reg_9_26_inst : DFFX1 port map( D => n841, CLK => n4879, Q => 
                           RAM_9_26_port, QN => n_2282);
   RAM_reg_9_25_inst : DFFX1 port map( D => n840, CLK => n4879, Q => 
                           RAM_9_25_port, QN => n_2283);
   RAM_reg_9_24_inst : DFFX1 port map( D => n839, CLK => n4879, Q => 
                           RAM_9_24_port, QN => n_2284);
   RAM_reg_9_23_inst : DFFX1 port map( D => n838, CLK => n4873, Q => 
                           RAM_9_23_port, QN => n_2285);
   RAM_reg_9_22_inst : DFFX1 port map( D => n837, CLK => n4873, Q => 
                           RAM_9_22_port, QN => n_2286);
   RAM_reg_9_21_inst : DFFX1 port map( D => n836, CLK => n4873, Q => 
                           RAM_9_21_port, QN => n_2287);
   RAM_reg_9_20_inst : DFFX1 port map( D => n835, CLK => n4873, Q => 
                           RAM_9_20_port, QN => n_2288);
   RAM_reg_9_19_inst : DFFX1 port map( D => n834, CLK => n4874, Q => 
                           RAM_9_19_port, QN => n_2289);
   RAM_reg_9_18_inst : DFFX1 port map( D => n833, CLK => n4874, Q => 
                           RAM_9_18_port, QN => n_2290);
   RAM_reg_9_17_inst : DFFX1 port map( D => n832, CLK => n4874, Q => 
                           RAM_9_17_port, QN => n_2291);
   RAM_reg_9_16_inst : DFFX1 port map( D => n831, CLK => n4874, Q => 
                           RAM_9_16_port, QN => n_2292);
   RAM_reg_9_15_inst : DFFX1 port map( D => n830, CLK => n4874, Q => 
                           RAM_9_15_port, QN => n_2293);
   RAM_reg_9_14_inst : DFFX1 port map( D => n829, CLK => n4874, Q => 
                           RAM_9_14_port, QN => n_2294);
   RAM_reg_9_13_inst : DFFX1 port map( D => n828, CLK => n4874, Q => 
                           RAM_9_13_port, QN => n_2295);
   RAM_reg_9_12_inst : DFFX1 port map( D => n827, CLK => n4874, Q => 
                           RAM_9_12_port, QN => n_2296);
   RAM_reg_9_11_inst : DFFX1 port map( D => n826, CLK => n4874, Q => 
                           RAM_9_11_port, QN => n_2297);
   RAM_reg_9_10_inst : DFFX1 port map( D => n825, CLK => n4874, Q => 
                           RAM_9_10_port, QN => n_2298);
   RAM_reg_9_9_inst : DFFX1 port map( D => n824, CLK => n4874, Q => 
                           RAM_9_9_port, QN => n_2299);
   RAM_reg_9_8_inst : DFFX1 port map( D => n823, CLK => n4874, Q => 
                           RAM_9_8_port, QN => n_2300);
   RAM_reg_9_7_inst : DFFX1 port map( D => n822, CLK => n4875, Q => 
                           RAM_9_7_port, QN => n_2301);
   RAM_reg_9_6_inst : DFFX1 port map( D => n821, CLK => n4875, Q => 
                           RAM_9_6_port, QN => n_2302);
   RAM_reg_9_5_inst : DFFX1 port map( D => n820, CLK => n4875, Q => 
                           RAM_9_5_port, QN => n_2303);
   RAM_reg_9_4_inst : DFFX1 port map( D => n819, CLK => n4875, Q => 
                           RAM_9_4_port, QN => n_2304);
   RAM_reg_9_3_inst : DFFX1 port map( D => n818, CLK => n4875, Q => 
                           RAM_9_3_port, QN => n_2305);
   RAM_reg_9_2_inst : DFFX1 port map( D => n817, CLK => n4875, Q => 
                           RAM_9_2_port, QN => n_2306);
   RAM_reg_9_1_inst : DFFX1 port map( D => n816, CLK => n4875, Q => 
                           RAM_9_1_port, QN => n_2307);
   RAM_reg_9_0_inst : DFFX1 port map( D => n815, CLK => n4875, Q => 
                           RAM_9_0_port, QN => n_2308);
   RAM_reg_10_127_inst : DFFX1 port map( D => n814, CLK => n4875, Q => 
                           RAM_10_127_port, QN => n_2309);
   RAM_reg_10_126_inst : DFFX1 port map( D => n813, CLK => n4875, Q => 
                           RAM_10_126_port, QN => n_2310);
   RAM_reg_10_125_inst : DFFX1 port map( D => n812, CLK => n4875, Q => 
                           RAM_10_125_port, QN => n_2311);
   RAM_reg_10_124_inst : DFFX1 port map( D => n811, CLK => n4875, Q => 
                           RAM_10_124_port, QN => n_2312);
   RAM_reg_10_123_inst : DFFX1 port map( D => n810, CLK => n4876, Q => 
                           RAM_10_123_port, QN => n_2313);
   RAM_reg_10_122_inst : DFFX1 port map( D => n809, CLK => n4876, Q => 
                           RAM_10_122_port, QN => n_2314);
   RAM_reg_10_121_inst : DFFX1 port map( D => n808, CLK => n4876, Q => 
                           RAM_10_121_port, QN => n_2315);
   RAM_reg_10_120_inst : DFFX1 port map( D => n807, CLK => n4876, Q => 
                           RAM_10_120_port, QN => n_2316);
   RAM_reg_10_119_inst : DFFX1 port map( D => n806, CLK => n4876, Q => 
                           RAM_10_119_port, QN => n_2317);
   RAM_reg_10_118_inst : DFFX1 port map( D => n805, CLK => n4876, Q => 
                           RAM_10_118_port, QN => n_2318);
   RAM_reg_10_117_inst : DFFX1 port map( D => n804, CLK => n4876, Q => 
                           RAM_10_117_port, QN => n_2319);
   RAM_reg_10_116_inst : DFFX1 port map( D => n803, CLK => n4876, Q => 
                           RAM_10_116_port, QN => n_2320);
   RAM_reg_10_115_inst : DFFX1 port map( D => n802, CLK => n4888, Q => 
                           RAM_10_115_port, QN => n_2321);
   RAM_reg_10_114_inst : DFFX1 port map( D => n801, CLK => n4888, Q => 
                           RAM_10_114_port, QN => n_2322);
   RAM_reg_10_113_inst : DFFX1 port map( D => n800, CLK => n4888, Q => 
                           RAM_10_113_port, QN => n_2323);
   RAM_reg_10_112_inst : DFFX1 port map( D => n799, CLK => n4888, Q => 
                           RAM_10_112_port, QN => n_2324);
   RAM_reg_10_111_inst : DFFX1 port map( D => n798, CLK => n4889, Q => 
                           RAM_10_111_port, QN => n_2325);
   RAM_reg_10_110_inst : DFFX1 port map( D => n797, CLK => n4889, Q => 
                           RAM_10_110_port, QN => n_2326);
   RAM_reg_10_109_inst : DFFX1 port map( D => n796, CLK => n4889, Q => 
                           RAM_10_109_port, QN => n_2327);
   RAM_reg_10_108_inst : DFFX1 port map( D => n795, CLK => n4889, Q => 
                           RAM_10_108_port, QN => n_2328);
   RAM_reg_10_107_inst : DFFX1 port map( D => n794, CLK => n4889, Q => 
                           RAM_10_107_port, QN => n_2329);
   RAM_reg_10_106_inst : DFFX1 port map( D => n793, CLK => n4889, Q => 
                           RAM_10_106_port, QN => n_2330);
   RAM_reg_10_105_inst : DFFX1 port map( D => n792, CLK => n4889, Q => 
                           RAM_10_105_port, QN => n_2331);
   RAM_reg_10_104_inst : DFFX1 port map( D => n791, CLK => n4889, Q => 
                           RAM_10_104_port, QN => n_2332);
   RAM_reg_10_103_inst : DFFX1 port map( D => n790, CLK => n4889, Q => 
                           RAM_10_103_port, QN => n_2333);
   RAM_reg_10_102_inst : DFFX1 port map( D => n789, CLK => n4889, Q => 
                           RAM_10_102_port, QN => n_2334);
   RAM_reg_10_101_inst : DFFX1 port map( D => n788, CLK => n4889, Q => 
                           RAM_10_101_port, QN => n_2335);
   RAM_reg_10_100_inst : DFFX1 port map( D => n787, CLK => n4889, Q => 
                           RAM_10_100_port, QN => n_2336);
   RAM_reg_10_99_inst : DFFX1 port map( D => n786, CLK => n4890, Q => 
                           RAM_10_99_port, QN => n_2337);
   RAM_reg_10_98_inst : DFFX1 port map( D => n785, CLK => n4890, Q => 
                           RAM_10_98_port, QN => n_2338);
   RAM_reg_10_97_inst : DFFX1 port map( D => n784, CLK => n4890, Q => 
                           RAM_10_97_port, QN => n_2339);
   RAM_reg_10_96_inst : DFFX1 port map( D => n783, CLK => n4890, Q => 
                           RAM_10_96_port, QN => n_2340);
   RAM_reg_10_95_inst : DFFX1 port map( D => n782, CLK => n4890, Q => 
                           RAM_10_95_port, QN => n_2341);
   RAM_reg_10_94_inst : DFFX1 port map( D => n781, CLK => n4890, Q => 
                           RAM_10_94_port, QN => n_2342);
   RAM_reg_10_93_inst : DFFX1 port map( D => n780, CLK => n4890, Q => 
                           RAM_10_93_port, QN => n_2343);
   RAM_reg_10_92_inst : DFFX1 port map( D => n779, CLK => n4890, Q => 
                           RAM_10_92_port, QN => n_2344);
   RAM_reg_10_91_inst : DFFX1 port map( D => n778, CLK => n4890, Q => 
                           RAM_10_91_port, QN => n_2345);
   RAM_reg_10_90_inst : DFFX1 port map( D => n777, CLK => n4890, Q => 
                           RAM_10_90_port, QN => n_2346);
   RAM_reg_10_89_inst : DFFX1 port map( D => n776, CLK => n4890, Q => 
                           RAM_10_89_port, QN => n_2347);
   RAM_reg_10_88_inst : DFFX1 port map( D => n775, CLK => n4890, Q => 
                           RAM_10_88_port, QN => n_2348);
   RAM_reg_10_87_inst : DFFX1 port map( D => n774, CLK => n4891, Q => 
                           RAM_10_87_port, QN => n_2349);
   RAM_reg_10_86_inst : DFFX1 port map( D => n773, CLK => n4891, Q => 
                           RAM_10_86_port, QN => n_2350);
   RAM_reg_10_85_inst : DFFX1 port map( D => n772, CLK => n4891, Q => 
                           RAM_10_85_port, QN => n_2351);
   RAM_reg_10_84_inst : DFFX1 port map( D => n771, CLK => n4891, Q => 
                           RAM_10_84_port, QN => n_2352);
   RAM_reg_10_83_inst : DFFX1 port map( D => n770, CLK => n4891, Q => 
                           RAM_10_83_port, QN => n_2353);
   RAM_reg_10_82_inst : DFFX1 port map( D => n769, CLK => n4891, Q => 
                           RAM_10_82_port, QN => n_2354);
   RAM_reg_10_81_inst : DFFX1 port map( D => n768, CLK => n4891, Q => 
                           RAM_10_81_port, QN => n_2355);
   RAM_reg_10_80_inst : DFFX1 port map( D => n767, CLK => n4891, Q => 
                           RAM_10_80_port, QN => n_2356);
   RAM_reg_10_79_inst : DFFX1 port map( D => n766, CLK => n4885, Q => 
                           RAM_10_79_port, QN => n_2357);
   RAM_reg_10_78_inst : DFFX1 port map( D => n765, CLK => n4885, Q => 
                           RAM_10_78_port, QN => n_2358);
   RAM_reg_10_77_inst : DFFX1 port map( D => n764, CLK => n4885, Q => 
                           RAM_10_77_port, QN => n_2359);
   RAM_reg_10_76_inst : DFFX1 port map( D => n763, CLK => n4885, Q => 
                           RAM_10_76_port, QN => n_2360);
   RAM_reg_10_75_inst : DFFX1 port map( D => n762, CLK => n4886, Q => 
                           RAM_10_75_port, QN => n_2361);
   RAM_reg_10_74_inst : DFFX1 port map( D => n761, CLK => n4886, Q => 
                           RAM_10_74_port, QN => n_2362);
   RAM_reg_10_73_inst : DFFX1 port map( D => n760, CLK => n4886, Q => 
                           RAM_10_73_port, QN => n_2363);
   RAM_reg_10_72_inst : DFFX1 port map( D => n759, CLK => n4886, Q => 
                           RAM_10_72_port, QN => n_2364);
   RAM_reg_10_71_inst : DFFX1 port map( D => n758, CLK => n4886, Q => 
                           RAM_10_71_port, QN => n_2365);
   RAM_reg_10_70_inst : DFFX1 port map( D => n757, CLK => n4886, Q => 
                           RAM_10_70_port, QN => n_2366);
   RAM_reg_10_69_inst : DFFX1 port map( D => n756, CLK => n4886, Q => 
                           RAM_10_69_port, QN => n_2367);
   RAM_reg_10_68_inst : DFFX1 port map( D => n755, CLK => n4886, Q => 
                           RAM_10_68_port, QN => n_2368);
   RAM_reg_10_67_inst : DFFX1 port map( D => n754, CLK => n4886, Q => 
                           RAM_10_67_port, QN => n_2369);
   RAM_reg_10_66_inst : DFFX1 port map( D => n753, CLK => n4886, Q => 
                           RAM_10_66_port, QN => n_2370);
   RAM_reg_10_65_inst : DFFX1 port map( D => n752, CLK => n4886, Q => 
                           RAM_10_65_port, QN => n_2371);
   RAM_reg_10_64_inst : DFFX1 port map( D => n751, CLK => n4886, Q => 
                           RAM_10_64_port, QN => n_2372);
   RAM_reg_10_63_inst : DFFX1 port map( D => n750, CLK => n4887, Q => 
                           RAM_10_63_port, QN => n_2373);
   RAM_reg_10_62_inst : DFFX1 port map( D => n749, CLK => n4887, Q => 
                           RAM_10_62_port, QN => n_2374);
   RAM_reg_10_61_inst : DFFX1 port map( D => n748, CLK => n4887, Q => 
                           RAM_10_61_port, QN => n_2375);
   RAM_reg_10_60_inst : DFFX1 port map( D => n747, CLK => n4887, Q => 
                           RAM_10_60_port, QN => n_2376);
   RAM_reg_10_59_inst : DFFX1 port map( D => n746, CLK => n4887, Q => 
                           RAM_10_59_port, QN => n_2377);
   RAM_reg_10_58_inst : DFFX1 port map( D => n745, CLK => n4887, Q => 
                           RAM_10_58_port, QN => n_2378);
   RAM_reg_10_57_inst : DFFX1 port map( D => n744, CLK => n4887, Q => 
                           RAM_10_57_port, QN => n_2379);
   RAM_reg_10_56_inst : DFFX1 port map( D => n743, CLK => n4887, Q => 
                           RAM_10_56_port, QN => n_2380);
   RAM_reg_10_55_inst : DFFX1 port map( D => n742, CLK => n4887, Q => 
                           RAM_10_55_port, QN => n_2381);
   RAM_reg_10_54_inst : DFFX1 port map( D => n741, CLK => n4887, Q => 
                           RAM_10_54_port, QN => n_2382);
   RAM_reg_10_53_inst : DFFX1 port map( D => n740, CLK => n4887, Q => 
                           RAM_10_53_port, QN => n_2383);
   RAM_reg_10_52_inst : DFFX1 port map( D => n739, CLK => n4887, Q => 
                           RAM_10_52_port, QN => n_2384);
   RAM_reg_10_51_inst : DFFX1 port map( D => n738, CLK => n4888, Q => 
                           RAM_10_51_port, QN => n_2385);
   RAM_reg_10_50_inst : DFFX1 port map( D => n737, CLK => n4888, Q => 
                           RAM_10_50_port, QN => n_2386);
   RAM_reg_10_49_inst : DFFX1 port map( D => n736, CLK => n4888, Q => 
                           RAM_10_49_port, QN => n_2387);
   RAM_reg_10_48_inst : DFFX1 port map( D => n735, CLK => n4888, Q => 
                           RAM_10_48_port, QN => n_2388);
   RAM_reg_10_47_inst : DFFX1 port map( D => n734, CLK => n4888, Q => 
                           RAM_10_47_port, QN => n_2389);
   RAM_reg_10_46_inst : DFFX1 port map( D => n733, CLK => n4888, Q => 
                           RAM_10_46_port, QN => n_2390);
   RAM_reg_10_45_inst : DFFX1 port map( D => n732, CLK => n4888, Q => 
                           RAM_10_45_port, QN => n_2391);
   RAM_reg_10_44_inst : DFFX1 port map( D => n731, CLK => n4888, Q => 
                           RAM_10_44_port, QN => n_2392);
   RAM_reg_10_43_inst : DFFX1 port map( D => n730, CLK => n4882, Q => 
                           RAM_10_43_port, QN => n_2393);
   RAM_reg_10_42_inst : DFFX1 port map( D => n729, CLK => n4882, Q => 
                           RAM_10_42_port, QN => n_2394);
   RAM_reg_10_41_inst : DFFX1 port map( D => n728, CLK => n4882, Q => 
                           RAM_10_41_port, QN => n_2395);
   RAM_reg_10_40_inst : DFFX1 port map( D => n727, CLK => n4882, Q => 
                           RAM_10_40_port, QN => n_2396);
   RAM_reg_10_39_inst : DFFX1 port map( D => n726, CLK => n4883, Q => 
                           RAM_10_39_port, QN => n_2397);
   RAM_reg_10_38_inst : DFFX1 port map( D => n725, CLK => n4883, Q => 
                           RAM_10_38_port, QN => n_2398);
   RAM_reg_10_37_inst : DFFX1 port map( D => n724, CLK => n4883, Q => 
                           RAM_10_37_port, QN => n_2399);
   RAM_reg_10_36_inst : DFFX1 port map( D => n723, CLK => n4883, Q => 
                           RAM_10_36_port, QN => n_2400);
   RAM_reg_10_35_inst : DFFX1 port map( D => n722, CLK => n4883, Q => 
                           RAM_10_35_port, QN => n_2401);
   RAM_reg_10_34_inst : DFFX1 port map( D => n721, CLK => n4883, Q => 
                           RAM_10_34_port, QN => n_2402);
   RAM_reg_10_33_inst : DFFX1 port map( D => n720, CLK => n4883, Q => 
                           RAM_10_33_port, QN => n_2403);
   RAM_reg_10_32_inst : DFFX1 port map( D => n719, CLK => n4883, Q => 
                           RAM_10_32_port, QN => n_2404);
   RAM_reg_10_31_inst : DFFX1 port map( D => n718, CLK => n4883, Q => 
                           RAM_10_31_port, QN => n_2405);
   RAM_reg_10_30_inst : DFFX1 port map( D => n717, CLK => n4883, Q => 
                           RAM_10_30_port, QN => n_2406);
   RAM_reg_10_29_inst : DFFX1 port map( D => n716, CLK => n4883, Q => 
                           RAM_10_29_port, QN => n_2407);
   RAM_reg_10_28_inst : DFFX1 port map( D => n715, CLK => n4883, Q => 
                           RAM_10_28_port, QN => n_2408);
   RAM_reg_10_27_inst : DFFX1 port map( D => n714, CLK => n4884, Q => 
                           RAM_10_27_port, QN => n_2409);
   RAM_reg_10_26_inst : DFFX1 port map( D => n713, CLK => n4884, Q => 
                           RAM_10_26_port, QN => n_2410);
   RAM_reg_10_25_inst : DFFX1 port map( D => n712, CLK => n4884, Q => 
                           RAM_10_25_port, QN => n_2411);
   RAM_reg_10_24_inst : DFFX1 port map( D => n711, CLK => n4884, Q => 
                           RAM_10_24_port, QN => n_2412);
   RAM_reg_10_23_inst : DFFX1 port map( D => n710, CLK => n4884, Q => 
                           RAM_10_23_port, QN => n_2413);
   RAM_reg_10_22_inst : DFFX1 port map( D => n709, CLK => n4884, Q => 
                           RAM_10_22_port, QN => n_2414);
   RAM_reg_10_21_inst : DFFX1 port map( D => n708, CLK => n4884, Q => 
                           RAM_10_21_port, QN => n_2415);
   RAM_reg_10_20_inst : DFFX1 port map( D => n707, CLK => n4884, Q => 
                           RAM_10_20_port, QN => n_2416);
   RAM_reg_10_19_inst : DFFX1 port map( D => n706, CLK => n4884, Q => 
                           RAM_10_19_port, QN => n_2417);
   RAM_reg_10_18_inst : DFFX1 port map( D => n705, CLK => n4884, Q => 
                           RAM_10_18_port, QN => n_2418);
   RAM_reg_10_17_inst : DFFX1 port map( D => n704, CLK => n4884, Q => 
                           RAM_10_17_port, QN => n_2419);
   RAM_reg_10_16_inst : DFFX1 port map( D => n703, CLK => n4884, Q => 
                           RAM_10_16_port, QN => n_2420);
   RAM_reg_10_15_inst : DFFX1 port map( D => n702, CLK => n4885, Q => 
                           RAM_10_15_port, QN => n_2421);
   RAM_reg_10_14_inst : DFFX1 port map( D => n701, CLK => n4885, Q => 
                           RAM_10_14_port, QN => n_2422);
   RAM_reg_10_13_inst : DFFX1 port map( D => n700, CLK => n4885, Q => 
                           RAM_10_13_port, QN => n_2423);
   RAM_reg_10_12_inst : DFFX1 port map( D => n699, CLK => n4885, Q => 
                           RAM_10_12_port, QN => n_2424);
   RAM_reg_10_11_inst : DFFX1 port map( D => n698, CLK => n4885, Q => 
                           RAM_10_11_port, QN => n_2425);
   RAM_reg_10_10_inst : DFFX1 port map( D => n697, CLK => n4885, Q => 
                           RAM_10_10_port, QN => n_2426);
   RAM_reg_10_9_inst : DFFX1 port map( D => n696, CLK => n4885, Q => 
                           RAM_10_9_port, QN => n_2427);
   RAM_reg_10_8_inst : DFFX1 port map( D => n695, CLK => n4885, Q => 
                           RAM_10_8_port, QN => n_2428);
   RAM_reg_10_7_inst : DFFX1 port map( D => n694, CLK => n4897, Q => 
                           RAM_10_7_port, QN => n_2429);
   RAM_reg_10_6_inst : DFFX1 port map( D => n693, CLK => n4897, Q => 
                           RAM_10_6_port, QN => n_2430);
   RAM_reg_10_5_inst : DFFX1 port map( D => n692, CLK => n4897, Q => 
                           RAM_10_5_port, QN => n_2431);
   RAM_reg_10_4_inst : DFFX1 port map( D => n691, CLK => n4897, Q => 
                           RAM_10_4_port, QN => n_2432);
   RAM_reg_10_3_inst : DFFX1 port map( D => n690, CLK => n4898, Q => 
                           RAM_10_3_port, QN => n_2433);
   RAM_reg_10_2_inst : DFFX1 port map( D => n689, CLK => n4898, Q => 
                           RAM_10_2_port, QN => n_2434);
   RAM_reg_10_1_inst : DFFX1 port map( D => n688, CLK => n4898, Q => 
                           RAM_10_1_port, QN => n_2435);
   RAM_reg_10_0_inst : DFFX1 port map( D => n687, CLK => n4898, Q => 
                           RAM_10_0_port, QN => n_2436);
   RAM_reg_11_127_inst : DFFX1 port map( D => n686, CLK => n4898, Q => 
                           RAM_11_127_port, QN => n_2437);
   RAM_reg_11_126_inst : DFFX1 port map( D => n685, CLK => n4898, Q => 
                           RAM_11_126_port, QN => n_2438);
   RAM_reg_11_125_inst : DFFX1 port map( D => n684, CLK => n4898, Q => 
                           RAM_11_125_port, QN => n_2439);
   RAM_reg_11_124_inst : DFFX1 port map( D => n683, CLK => n4898, Q => 
                           RAM_11_124_port, QN => n_2440);
   RAM_reg_11_123_inst : DFFX1 port map( D => n682, CLK => n4898, Q => 
                           RAM_11_123_port, QN => n_2441);
   RAM_reg_11_122_inst : DFFX1 port map( D => n681, CLK => n4898, Q => 
                           RAM_11_122_port, QN => n_2442);
   RAM_reg_11_121_inst : DFFX1 port map( D => n680, CLK => n4898, Q => 
                           RAM_11_121_port, QN => n_2443);
   RAM_reg_11_120_inst : DFFX1 port map( D => n679, CLK => n4898, Q => 
                           RAM_11_120_port, QN => n_2444);
   RAM_reg_11_119_inst : DFFX1 port map( D => n678, CLK => n4899, Q => 
                           RAM_11_119_port, QN => n_2445);
   RAM_reg_11_118_inst : DFFX1 port map( D => n677, CLK => n4899, Q => 
                           RAM_11_118_port, QN => n_2446);
   RAM_reg_11_117_inst : DFFX1 port map( D => n676, CLK => n4899, Q => 
                           RAM_11_117_port, QN => n_2447);
   RAM_reg_11_116_inst : DFFX1 port map( D => n675, CLK => n4899, Q => 
                           RAM_11_116_port, QN => n_2448);
   RAM_reg_11_115_inst : DFFX1 port map( D => n674, CLK => n4899, Q => 
                           RAM_11_115_port, QN => n_2449);
   RAM_reg_11_114_inst : DFFX1 port map( D => n673, CLK => n4899, Q => 
                           RAM_11_114_port, QN => n_2450);
   RAM_reg_11_113_inst : DFFX1 port map( D => n672, CLK => n4899, Q => 
                           RAM_11_113_port, QN => n_2451);
   RAM_reg_11_112_inst : DFFX1 port map( D => n671, CLK => n4899, Q => 
                           RAM_11_112_port, QN => n_2452);
   RAM_reg_11_111_inst : DFFX1 port map( D => n670, CLK => n4899, Q => 
                           RAM_11_111_port, QN => n_2453);
   RAM_reg_11_110_inst : DFFX1 port map( D => n669, CLK => n4899, Q => 
                           RAM_11_110_port, QN => n_2454);
   RAM_reg_11_109_inst : DFFX1 port map( D => n668, CLK => n4899, Q => 
                           RAM_11_109_port, QN => n_2455);
   RAM_reg_11_108_inst : DFFX1 port map( D => n667, CLK => n4899, Q => 
                           RAM_11_108_port, QN => n_2456);
   RAM_reg_11_107_inst : DFFX1 port map( D => n666, CLK => n4900, Q => 
                           RAM_11_107_port, QN => n_2457);
   RAM_reg_11_106_inst : DFFX1 port map( D => n665, CLK => n4900, Q => 
                           RAM_11_106_port, QN => n_2458);
   RAM_reg_11_105_inst : DFFX1 port map( D => n664, CLK => n4900, Q => 
                           RAM_11_105_port, QN => n_2459);
   RAM_reg_11_104_inst : DFFX1 port map( D => n663, CLK => n4900, Q => 
                           RAM_11_104_port, QN => n_2460);
   RAM_reg_11_103_inst : DFFX1 port map( D => n662, CLK => n4900, Q => 
                           RAM_11_103_port, QN => n_2461);
   RAM_reg_11_102_inst : DFFX1 port map( D => n661, CLK => n4900, Q => 
                           RAM_11_102_port, QN => n_2462);
   RAM_reg_11_101_inst : DFFX1 port map( D => n660, CLK => n4900, Q => 
                           RAM_11_101_port, QN => n_2463);
   RAM_reg_11_100_inst : DFFX1 port map( D => n659, CLK => n4900, Q => 
                           RAM_11_100_port, QN => n_2464);
   RAM_reg_11_99_inst : DFFX1 port map( D => n658, CLK => n4894, Q => 
                           RAM_11_99_port, QN => n_2465);
   RAM_reg_11_98_inst : DFFX1 port map( D => n657, CLK => n4894, Q => 
                           RAM_11_98_port, QN => n_2466);
   RAM_reg_11_97_inst : DFFX1 port map( D => n656, CLK => n4894, Q => 
                           RAM_11_97_port, QN => n_2467);
   RAM_reg_11_96_inst : DFFX1 port map( D => n655, CLK => n4894, Q => 
                           RAM_11_96_port, QN => n_2468);
   RAM_reg_11_95_inst : DFFX1 port map( D => n654, CLK => n4895, Q => 
                           RAM_11_95_port, QN => n_2469);
   RAM_reg_11_94_inst : DFFX1 port map( D => n653, CLK => n4895, Q => 
                           RAM_11_94_port, QN => n_2470);
   RAM_reg_11_93_inst : DFFX1 port map( D => n652, CLK => n4895, Q => 
                           RAM_11_93_port, QN => n_2471);
   RAM_reg_11_92_inst : DFFX1 port map( D => n651, CLK => n4895, Q => 
                           RAM_11_92_port, QN => n_2472);
   RAM_reg_11_91_inst : DFFX1 port map( D => n650, CLK => n4895, Q => 
                           RAM_11_91_port, QN => n_2473);
   RAM_reg_11_90_inst : DFFX1 port map( D => n649, CLK => n4895, Q => 
                           RAM_11_90_port, QN => n_2474);
   RAM_reg_11_89_inst : DFFX1 port map( D => n648, CLK => n4895, Q => 
                           RAM_11_89_port, QN => n_2475);
   RAM_reg_11_88_inst : DFFX1 port map( D => n647, CLK => n4895, Q => 
                           RAM_11_88_port, QN => n_2476);
   RAM_reg_11_87_inst : DFFX1 port map( D => n646, CLK => n4895, Q => 
                           RAM_11_87_port, QN => n_2477);
   RAM_reg_11_86_inst : DFFX1 port map( D => n645, CLK => n4895, Q => 
                           RAM_11_86_port, QN => n_2478);
   RAM_reg_11_85_inst : DFFX1 port map( D => n644, CLK => n4895, Q => 
                           RAM_11_85_port, QN => n_2479);
   RAM_reg_11_84_inst : DFFX1 port map( D => n643, CLK => n4895, Q => 
                           RAM_11_84_port, QN => n_2480);
   RAM_reg_11_83_inst : DFFX1 port map( D => n642, CLK => n4896, Q => 
                           RAM_11_83_port, QN => n_2481);
   RAM_reg_11_82_inst : DFFX1 port map( D => n641, CLK => n4896, Q => 
                           RAM_11_82_port, QN => n_2482);
   RAM_reg_11_81_inst : DFFX1 port map( D => n640, CLK => n4896, Q => 
                           RAM_11_81_port, QN => n_2483);
   RAM_reg_11_80_inst : DFFX1 port map( D => n639, CLK => n4896, Q => 
                           RAM_11_80_port, QN => n_2484);
   RAM_reg_11_79_inst : DFFX1 port map( D => n638, CLK => n4896, Q => 
                           RAM_11_79_port, QN => n_2485);
   RAM_reg_11_78_inst : DFFX1 port map( D => n637, CLK => n4896, Q => 
                           RAM_11_78_port, QN => n_2486);
   RAM_reg_11_77_inst : DFFX1 port map( D => n636, CLK => n4896, Q => 
                           RAM_11_77_port, QN => n_2487);
   RAM_reg_11_76_inst : DFFX1 port map( D => n635, CLK => n4896, Q => 
                           RAM_11_76_port, QN => n_2488);
   RAM_reg_11_75_inst : DFFX1 port map( D => n634, CLK => n4896, Q => 
                           RAM_11_75_port, QN => n_2489);
   RAM_reg_11_74_inst : DFFX1 port map( D => n633, CLK => n4896, Q => 
                           RAM_11_74_port, QN => n_2490);
   RAM_reg_11_73_inst : DFFX1 port map( D => n632, CLK => n4896, Q => 
                           RAM_11_73_port, QN => n_2491);
   RAM_reg_11_72_inst : DFFX1 port map( D => n631, CLK => n4896, Q => 
                           RAM_11_72_port, QN => n_2492);
   RAM_reg_11_71_inst : DFFX1 port map( D => n630, CLK => n4897, Q => 
                           RAM_11_71_port, QN => n_2493);
   RAM_reg_11_70_inst : DFFX1 port map( D => n629, CLK => n4897, Q => 
                           RAM_11_70_port, QN => n_2494);
   RAM_reg_11_69_inst : DFFX1 port map( D => n628, CLK => n4897, Q => 
                           RAM_11_69_port, QN => n_2495);
   RAM_reg_11_68_inst : DFFX1 port map( D => n627, CLK => n4897, Q => 
                           RAM_11_68_port, QN => n_2496);
   RAM_reg_11_67_inst : DFFX1 port map( D => n626, CLK => n4897, Q => 
                           RAM_11_67_port, QN => n_2497);
   RAM_reg_11_66_inst : DFFX1 port map( D => n625, CLK => n4897, Q => 
                           RAM_11_66_port, QN => n_2498);
   RAM_reg_11_65_inst : DFFX1 port map( D => n624, CLK => n4897, Q => 
                           RAM_11_65_port, QN => n_2499);
   RAM_reg_11_64_inst : DFFX1 port map( D => n623, CLK => n4897, Q => 
                           RAM_11_64_port, QN => n_2500);
   RAM_reg_11_63_inst : DFFX1 port map( D => n622, CLK => n4891, Q => 
                           RAM_11_63_port, QN => n_2501);
   RAM_reg_11_62_inst : DFFX1 port map( D => n621, CLK => n4891, Q => 
                           RAM_11_62_port, QN => n_2502);
   RAM_reg_11_61_inst : DFFX1 port map( D => n620, CLK => n4891, Q => 
                           RAM_11_61_port, QN => n_2503);
   RAM_reg_11_60_inst : DFFX1 port map( D => n619, CLK => n4891, Q => 
                           RAM_11_60_port, QN => n_2504);
   RAM_reg_11_59_inst : DFFX1 port map( D => n618, CLK => n4892, Q => 
                           RAM_11_59_port, QN => n_2505);
   RAM_reg_11_58_inst : DFFX1 port map( D => n617, CLK => n4892, Q => 
                           RAM_11_58_port, QN => n_2506);
   RAM_reg_11_57_inst : DFFX1 port map( D => n616, CLK => n4892, Q => 
                           RAM_11_57_port, QN => n_2507);
   RAM_reg_11_56_inst : DFFX1 port map( D => n615, CLK => n4892, Q => 
                           RAM_11_56_port, QN => n_2508);
   RAM_reg_11_55_inst : DFFX1 port map( D => n614, CLK => n4892, Q => 
                           RAM_11_55_port, QN => n_2509);
   RAM_reg_11_54_inst : DFFX1 port map( D => n613, CLK => n4892, Q => 
                           RAM_11_54_port, QN => n_2510);
   RAM_reg_11_53_inst : DFFX1 port map( D => n612, CLK => n4892, Q => 
                           RAM_11_53_port, QN => n_2511);
   RAM_reg_11_52_inst : DFFX1 port map( D => n611, CLK => n4892, Q => 
                           RAM_11_52_port, QN => n_2512);
   RAM_reg_11_51_inst : DFFX1 port map( D => n610, CLK => n4892, Q => 
                           RAM_11_51_port, QN => n_2513);
   RAM_reg_11_50_inst : DFFX1 port map( D => n609, CLK => n4892, Q => 
                           RAM_11_50_port, QN => n_2514);
   RAM_reg_11_49_inst : DFFX1 port map( D => n608, CLK => n4892, Q => 
                           RAM_11_49_port, QN => n_2515);
   RAM_reg_11_48_inst : DFFX1 port map( D => n607, CLK => n4892, Q => 
                           RAM_11_48_port, QN => n_2516);
   RAM_reg_11_47_inst : DFFX1 port map( D => n606, CLK => n4893, Q => 
                           RAM_11_47_port, QN => n_2517);
   RAM_reg_11_46_inst : DFFX1 port map( D => n605, CLK => n4893, Q => 
                           RAM_11_46_port, QN => n_2518);
   RAM_reg_11_45_inst : DFFX1 port map( D => n604, CLK => n4893, Q => 
                           RAM_11_45_port, QN => n_2519);
   RAM_reg_11_44_inst : DFFX1 port map( D => n603, CLK => n4893, Q => 
                           RAM_11_44_port, QN => n_2520);
   RAM_reg_11_43_inst : DFFX1 port map( D => n602, CLK => n4893, Q => 
                           RAM_11_43_port, QN => n_2521);
   RAM_reg_11_42_inst : DFFX1 port map( D => n601, CLK => n4893, Q => 
                           RAM_11_42_port, QN => n_2522);
   RAM_reg_11_41_inst : DFFX1 port map( D => n600, CLK => n4893, Q => 
                           RAM_11_41_port, QN => n_2523);
   RAM_reg_11_40_inst : DFFX1 port map( D => n599, CLK => n4893, Q => 
                           RAM_11_40_port, QN => n_2524);
   RAM_reg_11_39_inst : DFFX1 port map( D => n598, CLK => n4893, Q => 
                           RAM_11_39_port, QN => n_2525);
   RAM_reg_11_38_inst : DFFX1 port map( D => n597, CLK => n4893, Q => 
                           RAM_11_38_port, QN => n_2526);
   RAM_reg_11_37_inst : DFFX1 port map( D => n596, CLK => n4893, Q => 
                           RAM_11_37_port, QN => n_2527);
   RAM_reg_11_36_inst : DFFX1 port map( D => n595, CLK => n4893, Q => 
                           RAM_11_36_port, QN => n_2528);
   RAM_reg_11_35_inst : DFFX1 port map( D => n594, CLK => n4894, Q => 
                           RAM_11_35_port, QN => n_2529);
   RAM_reg_11_34_inst : DFFX1 port map( D => n593, CLK => n4894, Q => 
                           RAM_11_34_port, QN => n_2530);
   RAM_reg_11_33_inst : DFFX1 port map( D => n592, CLK => n4894, Q => 
                           RAM_11_33_port, QN => n_2531);
   RAM_reg_11_32_inst : DFFX1 port map( D => n591, CLK => n4894, Q => 
                           RAM_11_32_port, QN => n_2532);
   RAM_reg_11_31_inst : DFFX1 port map( D => n590, CLK => n4894, Q => 
                           RAM_11_31_port, QN => n_2533);
   RAM_reg_11_30_inst : DFFX1 port map( D => n589, CLK => n4894, Q => 
                           RAM_11_30_port, QN => n_2534);
   RAM_reg_11_29_inst : DFFX1 port map( D => n588, CLK => n4894, Q => 
                           RAM_11_29_port, QN => n_2535);
   RAM_reg_11_28_inst : DFFX1 port map( D => n587, CLK => n4894, Q => 
                           RAM_11_28_port, QN => n_2536);
   RAM_reg_11_27_inst : DFFX1 port map( D => n586, CLK => n4906, Q => 
                           RAM_11_27_port, QN => n_2537);
   RAM_reg_11_26_inst : DFFX1 port map( D => n585, CLK => n4906, Q => 
                           RAM_11_26_port, QN => n_2538);
   RAM_reg_11_25_inst : DFFX1 port map( D => n584, CLK => n4906, Q => 
                           RAM_11_25_port, QN => n_2539);
   RAM_reg_11_24_inst : DFFX1 port map( D => n583, CLK => n4906, Q => 
                           RAM_11_24_port, QN => n_2540);
   RAM_reg_11_23_inst : DFFX1 port map( D => n582, CLK => n4907, Q => 
                           RAM_11_23_port, QN => n_2541);
   RAM_reg_11_22_inst : DFFX1 port map( D => n581, CLK => n4907, Q => 
                           RAM_11_22_port, QN => n_2542);
   RAM_reg_11_21_inst : DFFX1 port map( D => n580, CLK => n4907, Q => 
                           RAM_11_21_port, QN => n_2543);
   RAM_reg_11_20_inst : DFFX1 port map( D => n579, CLK => n4907, Q => 
                           RAM_11_20_port, QN => n_2544);
   RAM_reg_11_19_inst : DFFX1 port map( D => n578, CLK => n4907, Q => 
                           RAM_11_19_port, QN => n_2545);
   RAM_reg_11_18_inst : DFFX1 port map( D => n577, CLK => n4907, Q => 
                           RAM_11_18_port, QN => n_2546);
   RAM_reg_11_17_inst : DFFX1 port map( D => n576, CLK => n4907, Q => 
                           RAM_11_17_port, QN => n_2547);
   RAM_reg_11_16_inst : DFFX1 port map( D => n575, CLK => n4907, Q => 
                           RAM_11_16_port, QN => n_2548);
   RAM_reg_11_15_inst : DFFX1 port map( D => n574, CLK => n4907, Q => 
                           RAM_11_15_port, QN => n_2549);
   RAM_reg_11_14_inst : DFFX1 port map( D => n573, CLK => n4907, Q => 
                           RAM_11_14_port, QN => n_2550);
   RAM_reg_11_13_inst : DFFX1 port map( D => n572, CLK => n4907, Q => 
                           RAM_11_13_port, QN => n_2551);
   RAM_reg_11_12_inst : DFFX1 port map( D => n571, CLK => n4907, Q => 
                           RAM_11_12_port, QN => n_2552);
   RAM_reg_11_11_inst : DFFX1 port map( D => n570, CLK => n4908, Q => 
                           RAM_11_11_port, QN => n_2553);
   RAM_reg_11_10_inst : DFFX1 port map( D => n569, CLK => n4908, Q => 
                           RAM_11_10_port, QN => n_2554);
   RAM_reg_11_9_inst : DFFX1 port map( D => n568, CLK => n4908, Q => 
                           RAM_11_9_port, QN => n_2555);
   RAM_reg_11_8_inst : DFFX1 port map( D => n567, CLK => n4908, Q => 
                           RAM_11_8_port, QN => n_2556);
   RAM_reg_11_7_inst : DFFX1 port map( D => n566, CLK => n4908, Q => 
                           RAM_11_7_port, QN => n_2557);
   RAM_reg_11_6_inst : DFFX1 port map( D => n565, CLK => n4908, Q => 
                           RAM_11_6_port, QN => n_2558);
   RAM_reg_11_5_inst : DFFX1 port map( D => n564, CLK => n4908, Q => 
                           RAM_11_5_port, QN => n_2559);
   RAM_reg_11_4_inst : DFFX1 port map( D => n563, CLK => n4908, Q => 
                           RAM_11_4_port, QN => n_2560);
   RAM_reg_11_3_inst : DFFX1 port map( D => n562, CLK => n4908, Q => 
                           RAM_11_3_port, QN => n_2561);
   RAM_reg_11_2_inst : DFFX1 port map( D => n561, CLK => n4908, Q => 
                           RAM_11_2_port, QN => n_2562);
   RAM_reg_11_1_inst : DFFX1 port map( D => n560, CLK => n4908, Q => 
                           RAM_11_1_port, QN => n_2563);
   RAM_reg_11_0_inst : DFFX1 port map( D => n559, CLK => n4908, Q => 
                           RAM_11_0_port, QN => n_2564);
   RAM_reg_12_127_inst : DFFX1 port map( D => n558, CLK => n4909, Q => 
                           RAM_12_127_port, QN => n_2565);
   RAM_reg_12_126_inst : DFFX1 port map( D => n557, CLK => n4909, Q => 
                           RAM_12_126_port, QN => n_2566);
   RAM_reg_12_125_inst : DFFX1 port map( D => n556, CLK => n4909, Q => 
                           RAM_12_125_port, QN => n_2567);
   RAM_reg_12_124_inst : DFFX1 port map( D => n555, CLK => n4909, Q => 
                           RAM_12_124_port, QN => n_2568);
   RAM_reg_12_123_inst : DFFX1 port map( D => n554, CLK => n4909, Q => 
                           RAM_12_123_port, QN => n_2569);
   RAM_reg_12_122_inst : DFFX1 port map( D => n553, CLK => n4909, Q => 
                           RAM_12_122_port, QN => n_2570);
   RAM_reg_12_121_inst : DFFX1 port map( D => n552, CLK => n4909, Q => 
                           RAM_12_121_port, QN => n_2571);
   RAM_reg_12_120_inst : DFFX1 port map( D => n551, CLK => n4909, Q => 
                           RAM_12_120_port, QN => n_2572);
   RAM_reg_12_119_inst : DFFX1 port map( D => n550, CLK => n4903, Q => 
                           RAM_12_119_port, QN => n_2573);
   RAM_reg_12_118_inst : DFFX1 port map( D => n549, CLK => n4903, Q => 
                           RAM_12_118_port, QN => n_2574);
   RAM_reg_12_117_inst : DFFX1 port map( D => n548, CLK => n4903, Q => 
                           RAM_12_117_port, QN => n_2575);
   RAM_reg_12_116_inst : DFFX1 port map( D => n547, CLK => n4903, Q => 
                           RAM_12_116_port, QN => n_2576);
   RAM_reg_12_115_inst : DFFX1 port map( D => n546, CLK => n4904, Q => 
                           RAM_12_115_port, QN => n_2577);
   RAM_reg_12_114_inst : DFFX1 port map( D => n545, CLK => n4904, Q => 
                           RAM_12_114_port, QN => n_2578);
   RAM_reg_12_113_inst : DFFX1 port map( D => n544, CLK => n4904, Q => 
                           RAM_12_113_port, QN => n_2579);
   RAM_reg_12_112_inst : DFFX1 port map( D => n543, CLK => n4904, Q => 
                           RAM_12_112_port, QN => n_2580);
   RAM_reg_12_111_inst : DFFX1 port map( D => n542, CLK => n4904, Q => 
                           RAM_12_111_port, QN => n_2581);
   RAM_reg_12_110_inst : DFFX1 port map( D => n541, CLK => n4904, Q => 
                           RAM_12_110_port, QN => n_2582);
   RAM_reg_12_109_inst : DFFX1 port map( D => n540, CLK => n4904, Q => 
                           RAM_12_109_port, QN => n_2583);
   RAM_reg_12_108_inst : DFFX1 port map( D => n539, CLK => n4904, Q => 
                           RAM_12_108_port, QN => n_2584);
   RAM_reg_12_107_inst : DFFX1 port map( D => n538, CLK => n4904, Q => 
                           RAM_12_107_port, QN => n_2585);
   RAM_reg_12_106_inst : DFFX1 port map( D => n537, CLK => n4904, Q => 
                           RAM_12_106_port, QN => n_2586);
   RAM_reg_12_105_inst : DFFX1 port map( D => n536, CLK => n4904, Q => 
                           RAM_12_105_port, QN => n_2587);
   RAM_reg_12_104_inst : DFFX1 port map( D => n535, CLK => n4904, Q => 
                           RAM_12_104_port, QN => n_2588);
   RAM_reg_12_103_inst : DFFX1 port map( D => n534, CLK => n4905, Q => 
                           RAM_12_103_port, QN => n_2589);
   RAM_reg_12_102_inst : DFFX1 port map( D => n533, CLK => n4905, Q => 
                           RAM_12_102_port, QN => n_2590);
   RAM_reg_12_101_inst : DFFX1 port map( D => n532, CLK => n4905, Q => 
                           RAM_12_101_port, QN => n_2591);
   RAM_reg_12_100_inst : DFFX1 port map( D => n531, CLK => n4905, Q => 
                           RAM_12_100_port, QN => n_2592);
   RAM_reg_12_99_inst : DFFX1 port map( D => n530, CLK => n4905, Q => 
                           RAM_12_99_port, QN => n_2593);
   RAM_reg_12_98_inst : DFFX1 port map( D => n529, CLK => n4905, Q => 
                           RAM_12_98_port, QN => n_2594);
   RAM_reg_12_97_inst : DFFX1 port map( D => n528, CLK => n4905, Q => 
                           RAM_12_97_port, QN => n_2595);
   RAM_reg_12_96_inst : DFFX1 port map( D => n527, CLK => n4905, Q => 
                           RAM_12_96_port, QN => n_2596);
   RAM_reg_12_95_inst : DFFX1 port map( D => n526, CLK => n4905, Q => 
                           RAM_12_95_port, QN => n_2597);
   RAM_reg_12_94_inst : DFFX1 port map( D => n525, CLK => n4905, Q => 
                           RAM_12_94_port, QN => n_2598);
   RAM_reg_12_93_inst : DFFX1 port map( D => n524, CLK => n4905, Q => 
                           RAM_12_93_port, QN => n_2599);
   RAM_reg_12_92_inst : DFFX1 port map( D => n523, CLK => n4905, Q => 
                           RAM_12_92_port, QN => n_2600);
   RAM_reg_12_91_inst : DFFX1 port map( D => n522, CLK => n4906, Q => 
                           RAM_12_91_port, QN => n_2601);
   RAM_reg_12_90_inst : DFFX1 port map( D => n521, CLK => n4906, Q => 
                           RAM_12_90_port, QN => n_2602);
   RAM_reg_12_89_inst : DFFX1 port map( D => n520, CLK => n4906, Q => 
                           RAM_12_89_port, QN => n_2603);
   RAM_reg_12_88_inst : DFFX1 port map( D => n519, CLK => n4906, Q => 
                           RAM_12_88_port, QN => n_2604);
   RAM_reg_12_87_inst : DFFX1 port map( D => n518, CLK => n4906, Q => 
                           RAM_12_87_port, QN => n_2605);
   RAM_reg_12_86_inst : DFFX1 port map( D => n517, CLK => n4906, Q => 
                           RAM_12_86_port, QN => n_2606);
   RAM_reg_12_85_inst : DFFX1 port map( D => n516, CLK => n4906, Q => 
                           RAM_12_85_port, QN => n_2607);
   RAM_reg_12_84_inst : DFFX1 port map( D => n515, CLK => n4906, Q => 
                           RAM_12_84_port, QN => n_2608);
   RAM_reg_12_83_inst : DFFX1 port map( D => n514, CLK => n4900, Q => 
                           RAM_12_83_port, QN => n_2609);
   RAM_reg_12_82_inst : DFFX1 port map( D => n513, CLK => n4900, Q => 
                           RAM_12_82_port, QN => n_2610);
   RAM_reg_12_81_inst : DFFX1 port map( D => n512, CLK => n4900, Q => 
                           RAM_12_81_port, QN => n_2611);
   RAM_reg_12_80_inst : DFFX1 port map( D => n511, CLK => n4900, Q => 
                           RAM_12_80_port, QN => n_2612);
   RAM_reg_12_79_inst : DFFX1 port map( D => n510, CLK => n4901, Q => 
                           RAM_12_79_port, QN => n_2613);
   RAM_reg_12_78_inst : DFFX1 port map( D => n509, CLK => n4901, Q => 
                           RAM_12_78_port, QN => n_2614);
   RAM_reg_12_77_inst : DFFX1 port map( D => n508, CLK => n4901, Q => 
                           RAM_12_77_port, QN => n_2615);
   RAM_reg_12_76_inst : DFFX1 port map( D => n507, CLK => n4901, Q => 
                           RAM_12_76_port, QN => n_2616);
   RAM_reg_12_75_inst : DFFX1 port map( D => n506, CLK => n4901, Q => 
                           RAM_12_75_port, QN => n_2617);
   RAM_reg_12_74_inst : DFFX1 port map( D => n505, CLK => n4901, Q => 
                           RAM_12_74_port, QN => n_2618);
   RAM_reg_12_73_inst : DFFX1 port map( D => n504, CLK => n4901, Q => 
                           RAM_12_73_port, QN => n_2619);
   RAM_reg_12_72_inst : DFFX1 port map( D => n503, CLK => n4901, Q => 
                           RAM_12_72_port, QN => n_2620);
   RAM_reg_12_71_inst : DFFX1 port map( D => n502, CLK => n4901, Q => 
                           RAM_12_71_port, QN => n_2621);
   RAM_reg_12_70_inst : DFFX1 port map( D => n501, CLK => n4901, Q => 
                           RAM_12_70_port, QN => n_2622);
   RAM_reg_12_69_inst : DFFX1 port map( D => n500, CLK => n4901, Q => 
                           RAM_12_69_port, QN => n_2623);
   RAM_reg_12_68_inst : DFFX1 port map( D => n499, CLK => n4901, Q => 
                           RAM_12_68_port, QN => n_2624);
   RAM_reg_12_67_inst : DFFX1 port map( D => n498, CLK => n4902, Q => 
                           RAM_12_67_port, QN => n_2625);
   RAM_reg_12_66_inst : DFFX1 port map( D => n497, CLK => n4902, Q => 
                           RAM_12_66_port, QN => n_2626);
   RAM_reg_12_65_inst : DFFX1 port map( D => n496, CLK => n4902, Q => 
                           RAM_12_65_port, QN => n_2627);
   RAM_reg_12_64_inst : DFFX1 port map( D => n495, CLK => n4902, Q => 
                           RAM_12_64_port, QN => n_2628);
   RAM_reg_12_63_inst : DFFX1 port map( D => n494, CLK => n4902, Q => 
                           RAM_12_63_port, QN => n_2629);
   RAM_reg_12_62_inst : DFFX1 port map( D => n493, CLK => n4902, Q => 
                           RAM_12_62_port, QN => n_2630);
   RAM_reg_12_61_inst : DFFX1 port map( D => n492, CLK => n4902, Q => 
                           RAM_12_61_port, QN => n_2631);
   RAM_reg_12_60_inst : DFFX1 port map( D => n491, CLK => n4902, Q => 
                           RAM_12_60_port, QN => n_2632);
   RAM_reg_12_59_inst : DFFX1 port map( D => n490, CLK => n4902, Q => 
                           RAM_12_59_port, QN => n_2633);
   RAM_reg_12_58_inst : DFFX1 port map( D => n489, CLK => n4902, Q => 
                           RAM_12_58_port, QN => n_2634);
   RAM_reg_12_57_inst : DFFX1 port map( D => n488, CLK => n4902, Q => 
                           RAM_12_57_port, QN => n_2635);
   RAM_reg_12_56_inst : DFFX1 port map( D => n487, CLK => n4902, Q => 
                           RAM_12_56_port, QN => n_2636);
   RAM_reg_12_55_inst : DFFX1 port map( D => n486, CLK => n4903, Q => 
                           RAM_12_55_port, QN => n_2637);
   RAM_reg_12_54_inst : DFFX1 port map( D => n485, CLK => n4903, Q => 
                           RAM_12_54_port, QN => n_2638);
   RAM_reg_12_53_inst : DFFX1 port map( D => n484, CLK => n4903, Q => 
                           RAM_12_53_port, QN => n_2639);
   RAM_reg_12_52_inst : DFFX1 port map( D => n483, CLK => n4903, Q => 
                           RAM_12_52_port, QN => n_2640);
   RAM_reg_12_51_inst : DFFX1 port map( D => n482, CLK => n4903, Q => 
                           RAM_12_51_port, QN => n_2641);
   RAM_reg_12_50_inst : DFFX1 port map( D => n481, CLK => n4903, Q => 
                           RAM_12_50_port, QN => n_2642);
   RAM_reg_12_49_inst : DFFX1 port map( D => n480, CLK => n4903, Q => 
                           RAM_12_49_port, QN => n_2643);
   RAM_reg_12_48_inst : DFFX1 port map( D => n479, CLK => n4903, Q => 
                           RAM_12_48_port, QN => n_2644);
   RAM_reg_12_47_inst : DFFX1 port map( D => n478, CLK => n4915, Q => 
                           RAM_12_47_port, QN => n_2645);
   RAM_reg_12_46_inst : DFFX1 port map( D => n477, CLK => n4915, Q => 
                           RAM_12_46_port, QN => n_2646);
   RAM_reg_12_45_inst : DFFX1 port map( D => n476, CLK => n4915, Q => 
                           RAM_12_45_port, QN => n_2647);
   RAM_reg_12_44_inst : DFFX1 port map( D => n475, CLK => n4915, Q => 
                           RAM_12_44_port, QN => n_2648);
   RAM_reg_12_43_inst : DFFX1 port map( D => n474, CLK => n4916, Q => 
                           RAM_12_43_port, QN => n_2649);
   RAM_reg_12_42_inst : DFFX1 port map( D => n473, CLK => n4916, Q => 
                           RAM_12_42_port, QN => n_2650);
   RAM_reg_12_41_inst : DFFX1 port map( D => n472, CLK => n4916, Q => 
                           RAM_12_41_port, QN => n_2651);
   RAM_reg_12_40_inst : DFFX1 port map( D => n471, CLK => n4916, Q => 
                           RAM_12_40_port, QN => n_2652);
   RAM_reg_12_39_inst : DFFX1 port map( D => n470, CLK => n4916, Q => 
                           RAM_12_39_port, QN => n_2653);
   RAM_reg_12_38_inst : DFFX1 port map( D => n469, CLK => n4916, Q => 
                           RAM_12_38_port, QN => n_2654);
   RAM_reg_12_37_inst : DFFX1 port map( D => n468, CLK => n4916, Q => 
                           RAM_12_37_port, QN => n_2655);
   RAM_reg_12_36_inst : DFFX1 port map( D => n467, CLK => n4916, Q => 
                           RAM_12_36_port, QN => n_2656);
   RAM_reg_12_35_inst : DFFX1 port map( D => n466, CLK => n4916, Q => 
                           RAM_12_35_port, QN => n_2657);
   RAM_reg_12_34_inst : DFFX1 port map( D => n465, CLK => n4916, Q => 
                           RAM_12_34_port, QN => n_2658);
   RAM_reg_12_33_inst : DFFX1 port map( D => n464, CLK => n4916, Q => 
                           RAM_12_33_port, QN => n_2659);
   RAM_reg_12_32_inst : DFFX1 port map( D => n463, CLK => n4916, Q => 
                           RAM_12_32_port, QN => n_2660);
   RAM_reg_12_31_inst : DFFX1 port map( D => n462, CLK => n4917, Q => 
                           RAM_12_31_port, QN => n_2661);
   RAM_reg_12_30_inst : DFFX1 port map( D => n461, CLK => n4917, Q => 
                           RAM_12_30_port, QN => n_2662);
   RAM_reg_12_29_inst : DFFX1 port map( D => n460, CLK => n4917, Q => 
                           RAM_12_29_port, QN => n_2663);
   RAM_reg_12_28_inst : DFFX1 port map( D => n459, CLK => n4917, Q => 
                           RAM_12_28_port, QN => n_2664);
   RAM_reg_12_27_inst : DFFX1 port map( D => n458, CLK => n4917, Q => 
                           RAM_12_27_port, QN => n_2665);
   RAM_reg_12_26_inst : DFFX1 port map( D => n457, CLK => n4917, Q => 
                           RAM_12_26_port, QN => n_2666);
   RAM_reg_12_25_inst : DFFX1 port map( D => n456, CLK => n4917, Q => 
                           RAM_12_25_port, QN => n_2667);
   RAM_reg_12_24_inst : DFFX1 port map( D => n455, CLK => n4917, Q => 
                           RAM_12_24_port, QN => n_2668);
   RAM_reg_12_23_inst : DFFX1 port map( D => n454, CLK => n4917, Q => 
                           RAM_12_23_port, QN => n_2669);
   RAM_reg_12_22_inst : DFFX1 port map( D => n453, CLK => n4917, Q => 
                           RAM_12_22_port, QN => n_2670);
   RAM_reg_12_21_inst : DFFX1 port map( D => n452, CLK => n4917, Q => 
                           RAM_12_21_port, QN => n_2671);
   RAM_reg_12_20_inst : DFFX1 port map( D => n451, CLK => n4917, Q => 
                           RAM_12_20_port, QN => n_2672);
   RAM_reg_12_19_inst : DFFX1 port map( D => n450, CLK => n4918, Q => 
                           RAM_12_19_port, QN => n_2673);
   RAM_reg_12_18_inst : DFFX1 port map( D => n449, CLK => n4918, Q => 
                           RAM_12_18_port, QN => n_2674);
   RAM_reg_12_17_inst : DFFX1 port map( D => n448, CLK => n4918, Q => 
                           RAM_12_17_port, QN => n_2675);
   RAM_reg_12_16_inst : DFFX1 port map( D => n447, CLK => n4918, Q => 
                           RAM_12_16_port, QN => n_2676);
   RAM_reg_12_15_inst : DFFX1 port map( D => n446, CLK => n4918, Q => 
                           RAM_12_15_port, QN => n_2677);
   RAM_reg_12_14_inst : DFFX1 port map( D => n445, CLK => n4918, Q => 
                           RAM_12_14_port, QN => n_2678);
   RAM_reg_12_13_inst : DFFX1 port map( D => n444, CLK => n4918, Q => 
                           RAM_12_13_port, QN => n_2679);
   RAM_reg_12_12_inst : DFFX1 port map( D => n443, CLK => n4918, Q => 
                           RAM_12_12_port, QN => n_2680);
   RAM_reg_12_11_inst : DFFX1 port map( D => n442, CLK => n4912, Q => 
                           RAM_12_11_port, QN => n_2681);
   RAM_reg_12_10_inst : DFFX1 port map( D => n441, CLK => n4912, Q => 
                           RAM_12_10_port, QN => n_2682);
   RAM_reg_12_9_inst : DFFX1 port map( D => n440, CLK => n4912, Q => 
                           RAM_12_9_port, QN => n_2683);
   RAM_reg_12_8_inst : DFFX1 port map( D => n439, CLK => n4912, Q => 
                           RAM_12_8_port, QN => n_2684);
   RAM_reg_12_7_inst : DFFX1 port map( D => n438, CLK => n4913, Q => 
                           RAM_12_7_port, QN => n_2685);
   RAM_reg_12_6_inst : DFFX1 port map( D => n437, CLK => n4913, Q => 
                           RAM_12_6_port, QN => n_2686);
   RAM_reg_12_5_inst : DFFX1 port map( D => n436, CLK => n4913, Q => 
                           RAM_12_5_port, QN => n_2687);
   RAM_reg_12_4_inst : DFFX1 port map( D => n435, CLK => n4913, Q => 
                           RAM_12_4_port, QN => n_2688);
   RAM_reg_12_3_inst : DFFX1 port map( D => n434, CLK => n4913, Q => 
                           RAM_12_3_port, QN => n_2689);
   RAM_reg_12_2_inst : DFFX1 port map( D => n433, CLK => n4913, Q => 
                           RAM_12_2_port, QN => n_2690);
   RAM_reg_12_1_inst : DFFX1 port map( D => n432, CLK => n4913, Q => 
                           RAM_12_1_port, QN => n_2691);
   RAM_reg_12_0_inst : DFFX1 port map( D => n431, CLK => n4913, Q => 
                           RAM_12_0_port, QN => n_2692);
   RAM_reg_13_127_inst : DFFX1 port map( D => n430, CLK => n4913, Q => 
                           RAM_13_127_port, QN => n_2693);
   RAM_reg_13_126_inst : DFFX1 port map( D => n429, CLK => n4913, Q => 
                           RAM_13_126_port, QN => n_2694);
   RAM_reg_13_125_inst : DFFX1 port map( D => n428, CLK => n4913, Q => 
                           RAM_13_125_port, QN => n_2695);
   RAM_reg_13_124_inst : DFFX1 port map( D => n427, CLK => n4913, Q => 
                           RAM_13_124_port, QN => n_2696);
   RAM_reg_13_123_inst : DFFX1 port map( D => n426, CLK => n4914, Q => 
                           RAM_13_123_port, QN => n_2697);
   RAM_reg_13_122_inst : DFFX1 port map( D => n425, CLK => n4914, Q => 
                           RAM_13_122_port, QN => n_2698);
   RAM_reg_13_121_inst : DFFX1 port map( D => n424, CLK => n4914, Q => 
                           RAM_13_121_port, QN => n_2699);
   RAM_reg_13_120_inst : DFFX1 port map( D => n423, CLK => n4914, Q => 
                           RAM_13_120_port, QN => n_2700);
   RAM_reg_13_119_inst : DFFX1 port map( D => n422, CLK => n4914, Q => 
                           RAM_13_119_port, QN => n_2701);
   RAM_reg_13_118_inst : DFFX1 port map( D => n421, CLK => n4914, Q => 
                           RAM_13_118_port, QN => n_2702);
   RAM_reg_13_117_inst : DFFX1 port map( D => n420, CLK => n4914, Q => 
                           RAM_13_117_port, QN => n_2703);
   RAM_reg_13_116_inst : DFFX1 port map( D => n419, CLK => n4914, Q => 
                           RAM_13_116_port, QN => n_2704);
   RAM_reg_13_115_inst : DFFX1 port map( D => n418, CLK => n4914, Q => 
                           RAM_13_115_port, QN => n_2705);
   RAM_reg_13_114_inst : DFFX1 port map( D => n417, CLK => n4914, Q => 
                           RAM_13_114_port, QN => n_2706);
   RAM_reg_13_113_inst : DFFX1 port map( D => n416, CLK => n4914, Q => 
                           RAM_13_113_port, QN => n_2707);
   RAM_reg_13_112_inst : DFFX1 port map( D => n415, CLK => n4914, Q => 
                           RAM_13_112_port, QN => n_2708);
   RAM_reg_13_111_inst : DFFX1 port map( D => n414, CLK => n4915, Q => 
                           RAM_13_111_port, QN => n_2709);
   RAM_reg_13_110_inst : DFFX1 port map( D => n413, CLK => n4915, Q => 
                           RAM_13_110_port, QN => n_2710);
   RAM_reg_13_109_inst : DFFX1 port map( D => n412, CLK => n4915, Q => 
                           RAM_13_109_port, QN => n_2711);
   RAM_reg_13_108_inst : DFFX1 port map( D => n411, CLK => n4915, Q => 
                           RAM_13_108_port, QN => n_2712);
   RAM_reg_13_107_inst : DFFX1 port map( D => n410, CLK => n4915, Q => 
                           RAM_13_107_port, QN => n_2713);
   RAM_reg_13_106_inst : DFFX1 port map( D => n409, CLK => n4915, Q => 
                           RAM_13_106_port, QN => n_2714);
   RAM_reg_13_105_inst : DFFX1 port map( D => n408, CLK => n4915, Q => 
                           RAM_13_105_port, QN => n_2715);
   RAM_reg_13_104_inst : DFFX1 port map( D => n407, CLK => n4915, Q => 
                           RAM_13_104_port, QN => n_2716);
   RAM_reg_13_103_inst : DFFX1 port map( D => n406, CLK => n4909, Q => 
                           RAM_13_103_port, QN => n_2717);
   RAM_reg_13_102_inst : DFFX1 port map( D => n405, CLK => n4909, Q => 
                           RAM_13_102_port, QN => n_2718);
   RAM_reg_13_101_inst : DFFX1 port map( D => n404, CLK => n4909, Q => 
                           RAM_13_101_port, QN => n_2719);
   RAM_reg_13_100_inst : DFFX1 port map( D => n403, CLK => n4909, Q => 
                           RAM_13_100_port, QN => n_2720);
   RAM_reg_13_99_inst : DFFX1 port map( D => n402, CLK => n4910, Q => 
                           RAM_13_99_port, QN => n_2721);
   RAM_reg_13_98_inst : DFFX1 port map( D => n401, CLK => n4910, Q => 
                           RAM_13_98_port, QN => n_2722);
   RAM_reg_13_97_inst : DFFX1 port map( D => n400, CLK => n4910, Q => 
                           RAM_13_97_port, QN => n_2723);
   RAM_reg_13_96_inst : DFFX1 port map( D => n399, CLK => n4910, Q => 
                           RAM_13_96_port, QN => n_2724);
   RAM_reg_13_95_inst : DFFX1 port map( D => n398, CLK => n4910, Q => 
                           RAM_13_95_port, QN => n_2725);
   RAM_reg_13_94_inst : DFFX1 port map( D => n397, CLK => n4910, Q => 
                           RAM_13_94_port, QN => n_2726);
   RAM_reg_13_93_inst : DFFX1 port map( D => n396, CLK => n4910, Q => 
                           RAM_13_93_port, QN => n_2727);
   RAM_reg_13_92_inst : DFFX1 port map( D => n395, CLK => n4910, Q => 
                           RAM_13_92_port, QN => n_2728);
   RAM_reg_13_91_inst : DFFX1 port map( D => n394, CLK => n4910, Q => 
                           RAM_13_91_port, QN => n_2729);
   RAM_reg_13_90_inst : DFFX1 port map( D => n393, CLK => n4910, Q => 
                           RAM_13_90_port, QN => n_2730);
   RAM_reg_13_89_inst : DFFX1 port map( D => n392, CLK => n4910, Q => 
                           RAM_13_89_port, QN => n_2731);
   RAM_reg_13_88_inst : DFFX1 port map( D => n391, CLK => n4910, Q => 
                           RAM_13_88_port, QN => n_2732);
   RAM_reg_13_87_inst : DFFX1 port map( D => n390, CLK => n4911, Q => 
                           RAM_13_87_port, QN => n_2733);
   RAM_reg_13_86_inst : DFFX1 port map( D => n389, CLK => n4911, Q => 
                           RAM_13_86_port, QN => n_2734);
   RAM_reg_13_85_inst : DFFX1 port map( D => n388, CLK => n4911, Q => 
                           RAM_13_85_port, QN => n_2735);
   RAM_reg_13_84_inst : DFFX1 port map( D => n387, CLK => n4911, Q => 
                           RAM_13_84_port, QN => n_2736);
   RAM_reg_13_83_inst : DFFX1 port map( D => n386, CLK => n4911, Q => 
                           RAM_13_83_port, QN => n_2737);
   RAM_reg_13_82_inst : DFFX1 port map( D => n385, CLK => n4911, Q => 
                           RAM_13_82_port, QN => n_2738);
   RAM_reg_13_81_inst : DFFX1 port map( D => n384, CLK => n4911, Q => 
                           RAM_13_81_port, QN => n_2739);
   RAM_reg_13_80_inst : DFFX1 port map( D => n383, CLK => n4911, Q => 
                           RAM_13_80_port, QN => n_2740);
   RAM_reg_13_79_inst : DFFX1 port map( D => n382, CLK => n4911, Q => 
                           RAM_13_79_port, QN => n_2741);
   RAM_reg_13_78_inst : DFFX1 port map( D => n381, CLK => n4911, Q => 
                           RAM_13_78_port, QN => n_2742);
   RAM_reg_13_77_inst : DFFX1 port map( D => n380, CLK => n4911, Q => 
                           RAM_13_77_port, QN => n_2743);
   RAM_reg_13_76_inst : DFFX1 port map( D => n379, CLK => n4911, Q => 
                           RAM_13_76_port, QN => n_2744);
   RAM_reg_13_75_inst : DFFX1 port map( D => n378, CLK => n4912, Q => 
                           RAM_13_75_port, QN => n_2745);
   RAM_reg_13_74_inst : DFFX1 port map( D => n377, CLK => n4912, Q => 
                           RAM_13_74_port, QN => n_2746);
   RAM_reg_13_73_inst : DFFX1 port map( D => n376, CLK => n4912, Q => 
                           RAM_13_73_port, QN => n_2747);
   RAM_reg_13_72_inst : DFFX1 port map( D => n375, CLK => n4912, Q => 
                           RAM_13_72_port, QN => n_2748);
   RAM_reg_13_71_inst : DFFX1 port map( D => n374, CLK => n4912, Q => 
                           RAM_13_71_port, QN => n_2749);
   RAM_reg_13_70_inst : DFFX1 port map( D => n373, CLK => n4912, Q => 
                           RAM_13_70_port, QN => n_2750);
   RAM_reg_13_69_inst : DFFX1 port map( D => n372, CLK => n4912, Q => 
                           RAM_13_69_port, QN => n_2751);
   RAM_reg_13_68_inst : DFFX1 port map( D => n371, CLK => n4912, Q => 
                           RAM_13_68_port, QN => n_2752);
   RAM_reg_13_67_inst : DFFX1 port map( D => n370, CLK => n4924, Q => 
                           RAM_13_67_port, QN => n_2753);
   RAM_reg_13_66_inst : DFFX1 port map( D => n369, CLK => n4924, Q => 
                           RAM_13_66_port, QN => n_2754);
   RAM_reg_13_65_inst : DFFX1 port map( D => n368, CLK => n4924, Q => 
                           RAM_13_65_port, QN => n_2755);
   RAM_reg_13_64_inst : DFFX1 port map( D => n367, CLK => n4924, Q => 
                           RAM_13_64_port, QN => n_2756);
   RAM_reg_13_63_inst : DFFX1 port map( D => n366, CLK => n4925, Q => 
                           RAM_13_63_port, QN => n_2757);
   RAM_reg_13_62_inst : DFFX1 port map( D => n365, CLK => n4925, Q => 
                           RAM_13_62_port, QN => n_2758);
   RAM_reg_13_61_inst : DFFX1 port map( D => n364, CLK => n4925, Q => 
                           RAM_13_61_port, QN => n_2759);
   RAM_reg_13_60_inst : DFFX1 port map( D => n363, CLK => n4925, Q => 
                           RAM_13_60_port, QN => n_2760);
   RAM_reg_13_59_inst : DFFX1 port map( D => n362, CLK => n4925, Q => 
                           RAM_13_59_port, QN => n_2761);
   RAM_reg_13_58_inst : DFFX1 port map( D => n361, CLK => n4925, Q => 
                           RAM_13_58_port, QN => n_2762);
   RAM_reg_13_57_inst : DFFX1 port map( D => n360, CLK => n4925, Q => 
                           RAM_13_57_port, QN => n_2763);
   RAM_reg_13_56_inst : DFFX1 port map( D => n359, CLK => n4925, Q => 
                           RAM_13_56_port, QN => n_2764);
   RAM_reg_13_55_inst : DFFX1 port map( D => n358, CLK => n4925, Q => 
                           RAM_13_55_port, QN => n_2765);
   RAM_reg_13_54_inst : DFFX1 port map( D => n357, CLK => n4925, Q => 
                           RAM_13_54_port, QN => n_2766);
   RAM_reg_13_53_inst : DFFX1 port map( D => n356, CLK => n4925, Q => 
                           RAM_13_53_port, QN => n_2767);
   RAM_reg_13_52_inst : DFFX1 port map( D => n355, CLK => n4925, Q => 
                           RAM_13_52_port, QN => n_2768);
   RAM_reg_13_51_inst : DFFX1 port map( D => n354, CLK => n4926, Q => 
                           RAM_13_51_port, QN => n_2769);
   RAM_reg_13_50_inst : DFFX1 port map( D => n353, CLK => n4926, Q => 
                           RAM_13_50_port, QN => n_2770);
   RAM_reg_13_49_inst : DFFX1 port map( D => n352, CLK => n4926, Q => 
                           RAM_13_49_port, QN => n_2771);
   RAM_reg_13_48_inst : DFFX1 port map( D => n351, CLK => n4926, Q => 
                           RAM_13_48_port, QN => n_2772);
   RAM_reg_13_47_inst : DFFX1 port map( D => n350, CLK => n4926, Q => 
                           RAM_13_47_port, QN => n_2773);
   RAM_reg_13_46_inst : DFFX1 port map( D => n349, CLK => n4926, Q => 
                           RAM_13_46_port, QN => n_2774);
   RAM_reg_13_45_inst : DFFX1 port map( D => n348, CLK => n4926, Q => 
                           RAM_13_45_port, QN => n_2775);
   RAM_reg_13_44_inst : DFFX1 port map( D => n347, CLK => n4926, Q => 
                           RAM_13_44_port, QN => n_2776);
   RAM_reg_13_43_inst : DFFX1 port map( D => n346, CLK => n4926, Q => 
                           RAM_13_43_port, QN => n_2777);
   RAM_reg_13_42_inst : DFFX1 port map( D => n345, CLK => n4926, Q => 
                           RAM_13_42_port, QN => n_2778);
   RAM_reg_13_41_inst : DFFX1 port map( D => n344, CLK => n4926, Q => 
                           RAM_13_41_port, QN => n_2779);
   RAM_reg_13_40_inst : DFFX1 port map( D => n343, CLK => n4926, Q => 
                           RAM_13_40_port, QN => n_2780);
   RAM_reg_13_39_inst : DFFX1 port map( D => n342, CLK => n4927, Q => 
                           RAM_13_39_port, QN => n_2781);
   RAM_reg_13_38_inst : DFFX1 port map( D => n341, CLK => n4927, Q => 
                           RAM_13_38_port, QN => n_2782);
   RAM_reg_13_37_inst : DFFX1 port map( D => n340, CLK => n4927, Q => 
                           RAM_13_37_port, QN => n_2783);
   RAM_reg_13_36_inst : DFFX1 port map( D => n339, CLK => n4927, Q => 
                           RAM_13_36_port, QN => n_2784);
   RAM_reg_13_35_inst : DFFX1 port map( D => n338, CLK => n4927, Q => 
                           RAM_13_35_port, QN => n_2785);
   RAM_reg_13_34_inst : DFFX1 port map( D => n337, CLK => n4927, Q => 
                           RAM_13_34_port, QN => n_2786);
   RAM_reg_13_33_inst : DFFX1 port map( D => n336, CLK => n4927, Q => 
                           RAM_13_33_port, QN => n_2787);
   RAM_reg_13_32_inst : DFFX1 port map( D => n335, CLK => n4927, Q => 
                           RAM_13_32_port, QN => n_2788);
   RAM_reg_13_31_inst : DFFX1 port map( D => n334, CLK => n4921, Q => 
                           RAM_13_31_port, QN => n_2789);
   RAM_reg_13_30_inst : DFFX1 port map( D => n333, CLK => n4921, Q => 
                           RAM_13_30_port, QN => n_2790);
   RAM_reg_13_29_inst : DFFX1 port map( D => n332, CLK => n4921, Q => 
                           RAM_13_29_port, QN => n_2791);
   RAM_reg_13_28_inst : DFFX1 port map( D => n331, CLK => n4921, Q => 
                           RAM_13_28_port, QN => n_2792);
   RAM_reg_13_27_inst : DFFX1 port map( D => n330, CLK => n4922, Q => 
                           RAM_13_27_port, QN => n_2793);
   RAM_reg_13_26_inst : DFFX1 port map( D => n329, CLK => n4922, Q => 
                           RAM_13_26_port, QN => n_2794);
   RAM_reg_13_25_inst : DFFX1 port map( D => n328, CLK => n4922, Q => 
                           RAM_13_25_port, QN => n_2795);
   RAM_reg_13_24_inst : DFFX1 port map( D => n327, CLK => n4922, Q => 
                           RAM_13_24_port, QN => n_2796);
   RAM_reg_13_23_inst : DFFX1 port map( D => n326, CLK => n4922, Q => 
                           RAM_13_23_port, QN => n_2797);
   RAM_reg_13_22_inst : DFFX1 port map( D => n325, CLK => n4922, Q => 
                           RAM_13_22_port, QN => n_2798);
   RAM_reg_13_21_inst : DFFX1 port map( D => n324, CLK => n4922, Q => 
                           RAM_13_21_port, QN => n_2799);
   RAM_reg_13_20_inst : DFFX1 port map( D => n323, CLK => n4922, Q => 
                           RAM_13_20_port, QN => n_2800);
   RAM_reg_13_19_inst : DFFX1 port map( D => n322, CLK => n4922, Q => 
                           RAM_13_19_port, QN => n_2801);
   RAM_reg_13_18_inst : DFFX1 port map( D => n321, CLK => n4922, Q => 
                           RAM_13_18_port, QN => n_2802);
   RAM_reg_13_17_inst : DFFX1 port map( D => n320, CLK => n4922, Q => 
                           RAM_13_17_port, QN => n_2803);
   RAM_reg_13_16_inst : DFFX1 port map( D => n319, CLK => n4922, Q => 
                           RAM_13_16_port, QN => n_2804);
   RAM_reg_13_15_inst : DFFX1 port map( D => n318, CLK => n4923, Q => 
                           RAM_13_15_port, QN => n_2805);
   RAM_reg_13_14_inst : DFFX1 port map( D => n317, CLK => n4923, Q => 
                           RAM_13_14_port, QN => n_2806);
   RAM_reg_13_13_inst : DFFX1 port map( D => n316, CLK => n4923, Q => 
                           RAM_13_13_port, QN => n_2807);
   RAM_reg_13_12_inst : DFFX1 port map( D => n315, CLK => n4923, Q => 
                           RAM_13_12_port, QN => n_2808);
   RAM_reg_13_11_inst : DFFX1 port map( D => n314, CLK => n4923, Q => 
                           RAM_13_11_port, QN => n_2809);
   RAM_reg_13_10_inst : DFFX1 port map( D => n313, CLK => n4923, Q => 
                           RAM_13_10_port, QN => n_2810);
   RAM_reg_13_9_inst : DFFX1 port map( D => n312, CLK => n4923, Q => 
                           RAM_13_9_port, QN => n_2811);
   RAM_reg_13_8_inst : DFFX1 port map( D => n311, CLK => n4923, Q => 
                           RAM_13_8_port, QN => n_2812);
   RAM_reg_13_7_inst : DFFX1 port map( D => n310, CLK => n4923, Q => 
                           RAM_13_7_port, QN => n_2813);
   RAM_reg_13_6_inst : DFFX1 port map( D => n309, CLK => n4923, Q => 
                           RAM_13_6_port, QN => n_2814);
   RAM_reg_13_5_inst : DFFX1 port map( D => n308, CLK => n4923, Q => 
                           RAM_13_5_port, QN => n_2815);
   RAM_reg_13_4_inst : DFFX1 port map( D => n307, CLK => n4923, Q => 
                           RAM_13_4_port, QN => n_2816);
   RAM_reg_13_3_inst : DFFX1 port map( D => n306, CLK => n4924, Q => 
                           RAM_13_3_port, QN => n_2817);
   RAM_reg_13_2_inst : DFFX1 port map( D => n305, CLK => n4924, Q => 
                           RAM_13_2_port, QN => n_2818);
   RAM_reg_13_1_inst : DFFX1 port map( D => n304, CLK => n4924, Q => 
                           RAM_13_1_port, QN => n_2819);
   RAM_reg_13_0_inst : DFFX1 port map( D => n303, CLK => n4924, Q => 
                           RAM_13_0_port, QN => n_2820);
   RAM_reg_14_127_inst : DFFX1 port map( D => n302, CLK => n4924, Q => 
                           RAM_14_127_port, QN => n_2821);
   RAM_reg_14_126_inst : DFFX1 port map( D => n301, CLK => n4924, Q => 
                           RAM_14_126_port, QN => n_2822);
   RAM_reg_14_125_inst : DFFX1 port map( D => n300, CLK => n4924, Q => 
                           RAM_14_125_port, QN => n_2823);
   RAM_reg_14_124_inst : DFFX1 port map( D => n299, CLK => n4924, Q => 
                           RAM_14_124_port, QN => n_2824);
   RAM_reg_14_123_inst : DFFX1 port map( D => n298, CLK => n4918, Q => 
                           RAM_14_123_port, QN => n_2825);
   RAM_reg_14_122_inst : DFFX1 port map( D => n297, CLK => n4918, Q => 
                           RAM_14_122_port, QN => n_2826);
   RAM_reg_14_121_inst : DFFX1 port map( D => n296, CLK => n4918, Q => 
                           RAM_14_121_port, QN => n_2827);
   RAM_reg_14_120_inst : DFFX1 port map( D => n295, CLK => n4918, Q => 
                           RAM_14_120_port, QN => n_2828);
   RAM_reg_14_119_inst : DFFX1 port map( D => n294, CLK => n4919, Q => 
                           RAM_14_119_port, QN => n_2829);
   RAM_reg_14_118_inst : DFFX1 port map( D => n293, CLK => n4919, Q => 
                           RAM_14_118_port, QN => n_2830);
   RAM_reg_14_117_inst : DFFX1 port map( D => n292, CLK => n4919, Q => 
                           RAM_14_117_port, QN => n_2831);
   RAM_reg_14_116_inst : DFFX1 port map( D => n291, CLK => n4919, Q => 
                           RAM_14_116_port, QN => n_2832);
   RAM_reg_14_115_inst : DFFX1 port map( D => n290, CLK => n4919, Q => 
                           RAM_14_115_port, QN => n_2833);
   RAM_reg_14_114_inst : DFFX1 port map( D => n289, CLK => n4919, Q => 
                           RAM_14_114_port, QN => n_2834);
   RAM_reg_14_113_inst : DFFX1 port map( D => n288, CLK => n4919, Q => 
                           RAM_14_113_port, QN => n_2835);
   RAM_reg_14_112_inst : DFFX1 port map( D => n287, CLK => n4919, Q => 
                           RAM_14_112_port, QN => n_2836);
   RAM_reg_14_111_inst : DFFX1 port map( D => n286, CLK => n4919, Q => 
                           RAM_14_111_port, QN => n_2837);
   RAM_reg_14_110_inst : DFFX1 port map( D => n285, CLK => n4919, Q => 
                           RAM_14_110_port, QN => n_2838);
   RAM_reg_14_109_inst : DFFX1 port map( D => n284, CLK => n4919, Q => 
                           RAM_14_109_port, QN => n_2839);
   RAM_reg_14_108_inst : DFFX1 port map( D => n283, CLK => n4919, Q => 
                           RAM_14_108_port, QN => n_2840);
   RAM_reg_14_107_inst : DFFX1 port map( D => n282, CLK => n4920, Q => 
                           RAM_14_107_port, QN => n_2841);
   RAM_reg_14_106_inst : DFFX1 port map( D => n281, CLK => n4920, Q => 
                           RAM_14_106_port, QN => n_2842);
   RAM_reg_14_105_inst : DFFX1 port map( D => n280, CLK => n4920, Q => 
                           RAM_14_105_port, QN => n_2843);
   RAM_reg_14_104_inst : DFFX1 port map( D => n279, CLK => n4920, Q => 
                           RAM_14_104_port, QN => n_2844);
   RAM_reg_14_103_inst : DFFX1 port map( D => n278, CLK => n4920, Q => 
                           RAM_14_103_port, QN => n_2845);
   RAM_reg_14_102_inst : DFFX1 port map( D => n277, CLK => n4920, Q => 
                           RAM_14_102_port, QN => n_2846);
   RAM_reg_14_101_inst : DFFX1 port map( D => n276, CLK => n4920, Q => 
                           RAM_14_101_port, QN => n_2847);
   RAM_reg_14_100_inst : DFFX1 port map( D => n275, CLK => n4920, Q => 
                           RAM_14_100_port, QN => n_2848);
   RAM_reg_14_99_inst : DFFX1 port map( D => n274, CLK => n4920, Q => 
                           RAM_14_99_port, QN => n_2849);
   RAM_reg_14_98_inst : DFFX1 port map( D => n273, CLK => n4920, Q => 
                           RAM_14_98_port, QN => n_2850);
   RAM_reg_14_97_inst : DFFX1 port map( D => n272, CLK => n4920, Q => 
                           RAM_14_97_port, QN => n_2851);
   RAM_reg_14_96_inst : DFFX1 port map( D => n271, CLK => n4920, Q => 
                           RAM_14_96_port, QN => n_2852);
   RAM_reg_14_95_inst : DFFX1 port map( D => n270, CLK => n4921, Q => 
                           RAM_14_95_port, QN => n_2853);
   RAM_reg_14_94_inst : DFFX1 port map( D => n269, CLK => n4921, Q => 
                           RAM_14_94_port, QN => n_2854);
   RAM_reg_14_93_inst : DFFX1 port map( D => n268, CLK => n4921, Q => 
                           RAM_14_93_port, QN => n_2855);
   RAM_reg_14_92_inst : DFFX1 port map( D => n267, CLK => n4921, Q => 
                           RAM_14_92_port, QN => n_2856);
   RAM_reg_14_91_inst : DFFX1 port map( D => n266, CLK => n4921, Q => 
                           RAM_14_91_port, QN => n_2857);
   RAM_reg_14_90_inst : DFFX1 port map( D => n265, CLK => n4921, Q => 
                           RAM_14_90_port, QN => n_2858);
   RAM_reg_14_89_inst : DFFX1 port map( D => n264, CLK => n4921, Q => 
                           RAM_14_89_port, QN => n_2859);
   RAM_reg_14_88_inst : DFFX1 port map( D => n263, CLK => n4921, Q => 
                           RAM_14_88_port, QN => n_2860);
   RAM_reg_14_87_inst : DFFX1 port map( D => n262, CLK => n4933, Q => 
                           RAM_14_87_port, QN => n_2861);
   RAM_reg_14_86_inst : DFFX1 port map( D => n261, CLK => n4933, Q => 
                           RAM_14_86_port, QN => n_2862);
   RAM_reg_14_85_inst : DFFX1 port map( D => n260, CLK => n4933, Q => 
                           RAM_14_85_port, QN => n_2863);
   RAM_reg_14_84_inst : DFFX1 port map( D => n259, CLK => n4933, Q => 
                           RAM_14_84_port, QN => n_2864);
   RAM_reg_14_83_inst : DFFX1 port map( D => n258, CLK => n4934, Q => 
                           RAM_14_83_port, QN => n_2865);
   RAM_reg_14_82_inst : DFFX1 port map( D => n257, CLK => n4934, Q => 
                           RAM_14_82_port, QN => n_2866);
   RAM_reg_14_81_inst : DFFX1 port map( D => n256, CLK => n4934, Q => 
                           RAM_14_81_port, QN => n_2867);
   RAM_reg_14_80_inst : DFFX1 port map( D => n255, CLK => n4934, Q => 
                           RAM_14_80_port, QN => n_2868);
   RAM_reg_14_79_inst : DFFX1 port map( D => n254, CLK => n4934, Q => 
                           RAM_14_79_port, QN => n_2869);
   RAM_reg_14_78_inst : DFFX1 port map( D => n253, CLK => n4934, Q => 
                           RAM_14_78_port, QN => n_2870);
   RAM_reg_14_77_inst : DFFX1 port map( D => n252, CLK => n4934, Q => 
                           RAM_14_77_port, QN => n_2871);
   RAM_reg_14_76_inst : DFFX1 port map( D => n251, CLK => n4934, Q => 
                           RAM_14_76_port, QN => n_2872);
   RAM_reg_14_75_inst : DFFX1 port map( D => n250, CLK => n4934, Q => 
                           RAM_14_75_port, QN => n_2873);
   RAM_reg_14_74_inst : DFFX1 port map( D => n249, CLK => n4934, Q => 
                           RAM_14_74_port, QN => n_2874);
   RAM_reg_14_73_inst : DFFX1 port map( D => n248, CLK => n4934, Q => 
                           RAM_14_73_port, QN => n_2875);
   RAM_reg_14_72_inst : DFFX1 port map( D => n247, CLK => n4934, Q => 
                           RAM_14_72_port, QN => n_2876);
   RAM_reg_14_71_inst : DFFX1 port map( D => n246, CLK => n4935, Q => 
                           RAM_14_71_port, QN => n_2877);
   RAM_reg_14_70_inst : DFFX1 port map( D => n245, CLK => n4935, Q => 
                           RAM_14_70_port, QN => n_2878);
   RAM_reg_14_69_inst : DFFX1 port map( D => n244, CLK => n4935, Q => 
                           RAM_14_69_port, QN => n_2879);
   RAM_reg_14_68_inst : DFFX1 port map( D => n243, CLK => n4935, Q => 
                           RAM_14_68_port, QN => n_2880);
   RAM_reg_14_67_inst : DFFX1 port map( D => n242, CLK => n4935, Q => 
                           RAM_14_67_port, QN => n_2881);
   RAM_reg_14_66_inst : DFFX1 port map( D => n241, CLK => n4935, Q => 
                           RAM_14_66_port, QN => n_2882);
   RAM_reg_14_65_inst : DFFX1 port map( D => n240, CLK => n4935, Q => 
                           RAM_14_65_port, QN => n_2883);
   RAM_reg_14_64_inst : DFFX1 port map( D => n239, CLK => n4935, Q => 
                           RAM_14_64_port, QN => n_2884);
   RAM_reg_14_63_inst : DFFX1 port map( D => n238, CLK => n4935, Q => 
                           RAM_14_63_port, QN => n_2885);
   RAM_reg_14_62_inst : DFFX1 port map( D => n237, CLK => n4935, Q => 
                           RAM_14_62_port, QN => n_2886);
   RAM_reg_14_61_inst : DFFX1 port map( D => n236, CLK => n4935, Q => 
                           RAM_14_61_port, QN => n_2887);
   RAM_reg_14_60_inst : DFFX1 port map( D => n235, CLK => n4935, Q => 
                           RAM_14_60_port, QN => n_2888);
   RAM_reg_14_59_inst : DFFX1 port map( D => n234, CLK => n4936, Q => 
                           RAM_14_59_port, QN => n_2889);
   RAM_reg_14_58_inst : DFFX1 port map( D => n233, CLK => n4936, Q => 
                           RAM_14_58_port, QN => n_2890);
   RAM_reg_14_57_inst : DFFX1 port map( D => n232, CLK => n4936, Q => 
                           RAM_14_57_port, QN => n_2891);
   RAM_reg_14_56_inst : DFFX1 port map( D => n231, CLK => n4936, Q => 
                           RAM_14_56_port, QN => n_2892);
   RAM_reg_14_55_inst : DFFX1 port map( D => n230, CLK => n4936, Q => 
                           RAM_14_55_port, QN => n_2893);
   RAM_reg_14_54_inst : DFFX1 port map( D => n229, CLK => n4936, Q => 
                           RAM_14_54_port, QN => n_2894);
   RAM_reg_14_53_inst : DFFX1 port map( D => n228, CLK => n4936, Q => 
                           RAM_14_53_port, QN => n_2895);
   RAM_reg_14_52_inst : DFFX1 port map( D => n227, CLK => n4936, Q => 
                           RAM_14_52_port, QN => n_2896);
   RAM_reg_14_51_inst : DFFX1 port map( D => n226, CLK => n4930, Q => 
                           RAM_14_51_port, QN => n_2897);
   RAM_reg_14_50_inst : DFFX1 port map( D => n225, CLK => n4930, Q => 
                           RAM_14_50_port, QN => n_2898);
   RAM_reg_14_49_inst : DFFX1 port map( D => n224, CLK => n4930, Q => 
                           RAM_14_49_port, QN => n_2899);
   RAM_reg_14_48_inst : DFFX1 port map( D => n223, CLK => n4930, Q => 
                           RAM_14_48_port, QN => n_2900);
   RAM_reg_14_47_inst : DFFX1 port map( D => n222, CLK => n4931, Q => 
                           RAM_14_47_port, QN => n_2901);
   RAM_reg_14_46_inst : DFFX1 port map( D => n221, CLK => n4931, Q => 
                           RAM_14_46_port, QN => n_2902);
   RAM_reg_14_45_inst : DFFX1 port map( D => n220, CLK => n4931, Q => 
                           RAM_14_45_port, QN => n_2903);
   RAM_reg_14_44_inst : DFFX1 port map( D => n219, CLK => n4931, Q => 
                           RAM_14_44_port, QN => n_2904);
   RAM_reg_14_43_inst : DFFX1 port map( D => n218, CLK => n4931, Q => 
                           RAM_14_43_port, QN => n_2905);
   RAM_reg_14_42_inst : DFFX1 port map( D => n217, CLK => n4931, Q => 
                           RAM_14_42_port, QN => n_2906);
   RAM_reg_14_41_inst : DFFX1 port map( D => n216, CLK => n4931, Q => 
                           RAM_14_41_port, QN => n_2907);
   RAM_reg_14_40_inst : DFFX1 port map( D => n215, CLK => n4931, Q => 
                           RAM_14_40_port, QN => n_2908);
   RAM_reg_14_39_inst : DFFX1 port map( D => n214, CLK => n4931, Q => 
                           RAM_14_39_port, QN => n_2909);
   RAM_reg_14_38_inst : DFFX1 port map( D => n213, CLK => n4931, Q => 
                           RAM_14_38_port, QN => n_2910);
   RAM_reg_14_37_inst : DFFX1 port map( D => n212, CLK => n4931, Q => 
                           RAM_14_37_port, QN => n_2911);
   RAM_reg_14_36_inst : DFFX1 port map( D => n211, CLK => n4931, Q => 
                           RAM_14_36_port, QN => n_2912);
   RAM_reg_14_35_inst : DFFX1 port map( D => n210, CLK => n4932, Q => 
                           RAM_14_35_port, QN => n_2913);
   RAM_reg_14_34_inst : DFFX1 port map( D => n209, CLK => n4932, Q => 
                           RAM_14_34_port, QN => n_2914);
   RAM_reg_14_33_inst : DFFX1 port map( D => n208, CLK => n4932, Q => 
                           RAM_14_33_port, QN => n_2915);
   RAM_reg_14_32_inst : DFFX1 port map( D => n207, CLK => n4932, Q => 
                           RAM_14_32_port, QN => n_2916);
   RAM_reg_14_31_inst : DFFX1 port map( D => n206, CLK => n4932, Q => 
                           RAM_14_31_port, QN => n_2917);
   RAM_reg_14_30_inst : DFFX1 port map( D => n205, CLK => n4932, Q => 
                           RAM_14_30_port, QN => n_2918);
   RAM_reg_14_29_inst : DFFX1 port map( D => n204, CLK => n4932, Q => 
                           RAM_14_29_port, QN => n_2919);
   RAM_reg_14_28_inst : DFFX1 port map( D => n203, CLK => n4932, Q => 
                           RAM_14_28_port, QN => n_2920);
   RAM_reg_14_27_inst : DFFX1 port map( D => n202, CLK => n4932, Q => 
                           RAM_14_27_port, QN => n_2921);
   RAM_reg_14_26_inst : DFFX1 port map( D => n201, CLK => n4932, Q => 
                           RAM_14_26_port, QN => n_2922);
   RAM_reg_14_25_inst : DFFX1 port map( D => n200, CLK => n4932, Q => 
                           RAM_14_25_port, QN => n_2923);
   RAM_reg_14_24_inst : DFFX1 port map( D => n199, CLK => n4932, Q => 
                           RAM_14_24_port, QN => n_2924);
   RAM_reg_14_23_inst : DFFX1 port map( D => n198, CLK => n4933, Q => 
                           RAM_14_23_port, QN => n_2925);
   RAM_reg_14_22_inst : DFFX1 port map( D => n197, CLK => n4933, Q => 
                           RAM_14_22_port, QN => n_2926);
   RAM_reg_14_21_inst : DFFX1 port map( D => n196, CLK => n4933, Q => 
                           RAM_14_21_port, QN => n_2927);
   RAM_reg_14_20_inst : DFFX1 port map( D => n195, CLK => n4933, Q => 
                           RAM_14_20_port, QN => n_2928);
   RAM_reg_14_19_inst : DFFX1 port map( D => n194, CLK => n4933, Q => 
                           RAM_14_19_port, QN => n_2929);
   RAM_reg_14_18_inst : DFFX1 port map( D => n193, CLK => n4933, Q => 
                           RAM_14_18_port, QN => n_2930);
   RAM_reg_14_17_inst : DFFX1 port map( D => n192, CLK => n4933, Q => 
                           RAM_14_17_port, QN => n_2931);
   RAM_reg_14_16_inst : DFFX1 port map( D => n191, CLK => n4933, Q => 
                           RAM_14_16_port, QN => n_2932);
   RAM_reg_14_15_inst : DFFX1 port map( D => n190, CLK => n4927, Q => 
                           RAM_14_15_port, QN => n_2933);
   RAM_reg_14_14_inst : DFFX1 port map( D => n189, CLK => n4927, Q => 
                           RAM_14_14_port, QN => n_2934);
   RAM_reg_14_13_inst : DFFX1 port map( D => n188, CLK => n4927, Q => 
                           RAM_14_13_port, QN => n_2935);
   RAM_reg_14_12_inst : DFFX1 port map( D => n187, CLK => n4927, Q => 
                           RAM_14_12_port, QN => n_2936);
   RAM_reg_14_11_inst : DFFX1 port map( D => n186, CLK => n4928, Q => 
                           RAM_14_11_port, QN => n_2937);
   RAM_reg_14_10_inst : DFFX1 port map( D => n185, CLK => n4928, Q => 
                           RAM_14_10_port, QN => n_2938);
   RAM_reg_14_9_inst : DFFX1 port map( D => n184, CLK => n4928, Q => 
                           RAM_14_9_port, QN => n_2939);
   RAM_reg_14_8_inst : DFFX1 port map( D => n183, CLK => n4928, Q => 
                           RAM_14_8_port, QN => n_2940);
   RAM_reg_14_7_inst : DFFX1 port map( D => n182, CLK => n4928, Q => 
                           RAM_14_7_port, QN => n_2941);
   RAM_reg_14_6_inst : DFFX1 port map( D => n181, CLK => n4928, Q => 
                           RAM_14_6_port, QN => n_2942);
   RAM_reg_14_5_inst : DFFX1 port map( D => n180, CLK => n4928, Q => 
                           RAM_14_5_port, QN => n_2943);
   RAM_reg_14_4_inst : DFFX1 port map( D => n179, CLK => n4928, Q => 
                           RAM_14_4_port, QN => n_2944);
   RAM_reg_14_3_inst : DFFX1 port map( D => n178, CLK => n4928, Q => 
                           RAM_14_3_port, QN => n_2945);
   RAM_reg_14_2_inst : DFFX1 port map( D => n177, CLK => n4928, Q => 
                           RAM_14_2_port, QN => n_2946);
   RAM_reg_14_1_inst : DFFX1 port map( D => n176, CLK => n4928, Q => 
                           RAM_14_1_port, QN => n_2947);
   RAM_reg_14_0_inst : DFFX1 port map( D => n175, CLK => n4928, Q => 
                           RAM_14_0_port, QN => n_2948);
   RAM_reg_15_127_inst : DFFX1 port map( D => n174, CLK => n4929, Q => 
                           RAM_15_127_port, QN => n_2949);
   RAM_reg_15_126_inst : DFFX1 port map( D => n173, CLK => n4929, Q => 
                           RAM_15_126_port, QN => n_2950);
   RAM_reg_15_125_inst : DFFX1 port map( D => n172, CLK => n4929, Q => 
                           RAM_15_125_port, QN => n_2951);
   RAM_reg_15_124_inst : DFFX1 port map( D => n171, CLK => n4929, Q => 
                           RAM_15_124_port, QN => n_2952);
   RAM_reg_15_123_inst : DFFX1 port map( D => n170, CLK => n4929, Q => 
                           RAM_15_123_port, QN => n_2953);
   RAM_reg_15_122_inst : DFFX1 port map( D => n169, CLK => n4929, Q => 
                           RAM_15_122_port, QN => n_2954);
   RAM_reg_15_121_inst : DFFX1 port map( D => n168, CLK => n4929, Q => 
                           RAM_15_121_port, QN => n_2955);
   RAM_reg_15_120_inst : DFFX1 port map( D => n167, CLK => n4929, Q => 
                           RAM_15_120_port, QN => n_2956);
   RAM_reg_15_119_inst : DFFX1 port map( D => n166, CLK => n4929, Q => 
                           RAM_15_119_port, QN => n_2957);
   RAM_reg_15_118_inst : DFFX1 port map( D => n165, CLK => n4929, Q => 
                           RAM_15_118_port, QN => n_2958);
   RAM_reg_15_117_inst : DFFX1 port map( D => n164, CLK => n4929, Q => 
                           RAM_15_117_port, QN => n_2959);
   RAM_reg_15_116_inst : DFFX1 port map( D => n163, CLK => n4929, Q => 
                           RAM_15_116_port, QN => n_2960);
   RAM_reg_15_115_inst : DFFX1 port map( D => n162, CLK => n4930, Q => 
                           RAM_15_115_port, QN => n_2961);
   RAM_reg_15_114_inst : DFFX1 port map( D => n161, CLK => n4930, Q => 
                           RAM_15_114_port, QN => n_2962);
   RAM_reg_15_113_inst : DFFX1 port map( D => n160, CLK => n4930, Q => 
                           RAM_15_113_port, QN => n_2963);
   RAM_reg_15_112_inst : DFFX1 port map( D => n159, CLK => n4930, Q => 
                           RAM_15_112_port, QN => n_2964);
   RAM_reg_15_111_inst : DFFX1 port map( D => n158, CLK => n4930, Q => 
                           RAM_15_111_port, QN => n_2965);
   RAM_reg_15_110_inst : DFFX1 port map( D => n157, CLK => n4930, Q => 
                           RAM_15_110_port, QN => n_2966);
   RAM_reg_15_109_inst : DFFX1 port map( D => n156, CLK => n4930, Q => 
                           RAM_15_109_port, QN => n_2967);
   RAM_reg_15_108_inst : DFFX1 port map( D => n155, CLK => n4930, Q => 
                           RAM_15_108_port, QN => n_2968);
   RAM_reg_15_107_inst : DFFX1 port map( D => n154, CLK => n4942, Q => 
                           RAM_15_107_port, QN => n_2969);
   RAM_reg_15_106_inst : DFFX1 port map( D => n153, CLK => n4942, Q => 
                           RAM_15_106_port, QN => n_2970);
   RAM_reg_15_105_inst : DFFX1 port map( D => n152, CLK => n4942, Q => 
                           RAM_15_105_port, QN => n_2971);
   RAM_reg_15_104_inst : DFFX1 port map( D => n151, CLK => n4942, Q => 
                           RAM_15_104_port, QN => n_2972);
   RAM_reg_15_103_inst : DFFX1 port map( D => n150, CLK => n4943, Q => 
                           RAM_15_103_port, QN => n_2973);
   RAM_reg_15_102_inst : DFFX1 port map( D => n149, CLK => n4943, Q => 
                           RAM_15_102_port, QN => n_2974);
   RAM_reg_15_101_inst : DFFX1 port map( D => n148, CLK => n4943, Q => 
                           RAM_15_101_port, QN => n_2975);
   RAM_reg_15_100_inst : DFFX1 port map( D => n147, CLK => n4943, Q => 
                           RAM_15_100_port, QN => n_2976);
   RAM_reg_15_99_inst : DFFX1 port map( D => n146, CLK => n4943, Q => 
                           RAM_15_99_port, QN => n_2977);
   RAM_reg_15_98_inst : DFFX1 port map( D => n145, CLK => n4943, Q => 
                           RAM_15_98_port, QN => n_2978);
   RAM_reg_15_97_inst : DFFX1 port map( D => n144, CLK => n4943, Q => 
                           RAM_15_97_port, QN => n_2979);
   RAM_reg_15_96_inst : DFFX1 port map( D => n143, CLK => n4943, Q => 
                           RAM_15_96_port, QN => n_2980);
   RAM_reg_15_95_inst : DFFX1 port map( D => n142, CLK => n4943, Q => 
                           RAM_15_95_port, QN => n_2981);
   RAM_reg_15_94_inst : DFFX1 port map( D => n141, CLK => n4943, Q => 
                           RAM_15_94_port, QN => n_2982);
   RAM_reg_15_93_inst : DFFX1 port map( D => n140, CLK => n4943, Q => 
                           RAM_15_93_port, QN => n_2983);
   RAM_reg_15_92_inst : DFFX1 port map( D => n139, CLK => n4943, Q => 
                           RAM_15_92_port, QN => n_2984);
   RAM_reg_15_91_inst : DFFX1 port map( D => n138, CLK => n4944, Q => 
                           RAM_15_91_port, QN => n_2985);
   RAM_reg_15_90_inst : DFFX1 port map( D => n137, CLK => n4944, Q => 
                           RAM_15_90_port, QN => n_2986);
   RAM_reg_15_89_inst : DFFX1 port map( D => n136, CLK => n4944, Q => 
                           RAM_15_89_port, QN => n_2987);
   RAM_reg_15_88_inst : DFFX1 port map( D => n135, CLK => n4944, Q => 
                           RAM_15_88_port, QN => n_2988);
   RAM_reg_15_87_inst : DFFX1 port map( D => n134, CLK => n4944, Q => 
                           RAM_15_87_port, QN => n_2989);
   RAM_reg_15_86_inst : DFFX1 port map( D => n133, CLK => n4944, Q => 
                           RAM_15_86_port, QN => n_2990);
   RAM_reg_15_85_inst : DFFX1 port map( D => n132, CLK => n4944, Q => 
                           RAM_15_85_port, QN => n_2991);
   RAM_reg_15_84_inst : DFFX1 port map( D => n131, CLK => n4944, Q => 
                           RAM_15_84_port, QN => n_2992);
   RAM_reg_15_83_inst : DFFX1 port map( D => n130, CLK => n4944, Q => 
                           RAM_15_83_port, QN => n_2993);
   RAM_reg_15_82_inst : DFFX1 port map( D => n129, CLK => n4944, Q => 
                           RAM_15_82_port, QN => n_2994);
   RAM_reg_15_81_inst : DFFX1 port map( D => n128, CLK => n4944, Q => 
                           RAM_15_81_port, QN => n_2995);
   RAM_reg_15_80_inst : DFFX1 port map( D => n127, CLK => n4944, Q => 
                           RAM_15_80_port, QN => n_2996);
   RAM_reg_15_79_inst : DFFX1 port map( D => n126, CLK => n4945, Q => 
                           RAM_15_79_port, QN => n_2997);
   RAM_reg_15_78_inst : DFFX1 port map( D => n125, CLK => n4945, Q => 
                           RAM_15_78_port, QN => n_2998);
   RAM_reg_15_77_inst : DFFX1 port map( D => n124, CLK => n4945, Q => 
                           RAM_15_77_port, QN => n_2999);
   RAM_reg_15_76_inst : DFFX1 port map( D => n123, CLK => n4945, Q => 
                           RAM_15_76_port, QN => n_3000);
   RAM_reg_15_75_inst : DFFX1 port map( D => n122, CLK => n4945, Q => 
                           RAM_15_75_port, QN => n_3001);
   RAM_reg_15_74_inst : DFFX1 port map( D => n121, CLK => n4945, Q => 
                           RAM_15_74_port, QN => n_3002);
   RAM_reg_15_73_inst : DFFX1 port map( D => n120, CLK => n4945, Q => 
                           RAM_15_73_port, QN => n_3003);
   RAM_reg_15_72_inst : DFFX1 port map( D => n119, CLK => n4945, Q => 
                           RAM_15_72_port, QN => n_3004);
   RAM_reg_15_71_inst : DFFX1 port map( D => n118, CLK => n4939, Q => 
                           RAM_15_71_port, QN => n_3005);
   RAM_reg_15_70_inst : DFFX1 port map( D => n117, CLK => n4939, Q => 
                           RAM_15_70_port, QN => n_3006);
   RAM_reg_15_69_inst : DFFX1 port map( D => n116, CLK => n4939, Q => 
                           RAM_15_69_port, QN => n_3007);
   RAM_reg_15_68_inst : DFFX1 port map( D => n115, CLK => n4939, Q => 
                           RAM_15_68_port, QN => n_3008);
   RAM_reg_15_67_inst : DFFX1 port map( D => n114, CLK => n4940, Q => 
                           RAM_15_67_port, QN => n_3009);
   RAM_reg_15_66_inst : DFFX1 port map( D => n113, CLK => n4940, Q => 
                           RAM_15_66_port, QN => n_3010);
   RAM_reg_15_65_inst : DFFX1 port map( D => n112, CLK => n4940, Q => 
                           RAM_15_65_port, QN => n_3011);
   RAM_reg_15_64_inst : DFFX1 port map( D => n111, CLK => n4940, Q => 
                           RAM_15_64_port, QN => n_3012);
   RAM_reg_15_63_inst : DFFX1 port map( D => n110, CLK => n4940, Q => 
                           RAM_15_63_port, QN => n_3013);
   RAM_reg_15_62_inst : DFFX1 port map( D => n109, CLK => n4940, Q => 
                           RAM_15_62_port, QN => n_3014);
   RAM_reg_15_61_inst : DFFX1 port map( D => n108, CLK => n4940, Q => 
                           RAM_15_61_port, QN => n_3015);
   RAM_reg_15_60_inst : DFFX1 port map( D => n107, CLK => n4940, Q => 
                           RAM_15_60_port, QN => n_3016);
   RAM_reg_15_59_inst : DFFX1 port map( D => n106, CLK => n4940, Q => 
                           RAM_15_59_port, QN => n_3017);
   RAM_reg_15_58_inst : DFFX1 port map( D => n105, CLK => n4940, Q => 
                           RAM_15_58_port, QN => n_3018);
   RAM_reg_15_57_inst : DFFX1 port map( D => n104, CLK => n4940, Q => 
                           RAM_15_57_port, QN => n_3019);
   RAM_reg_15_56_inst : DFFX1 port map( D => n103, CLK => n4940, Q => 
                           RAM_15_56_port, QN => n_3020);
   RAM_reg_15_55_inst : DFFX1 port map( D => n102, CLK => n4941, Q => 
                           RAM_15_55_port, QN => n_3021);
   RAM_reg_15_54_inst : DFFX1 port map( D => n101, CLK => n4941, Q => 
                           RAM_15_54_port, QN => n_3022);
   RAM_reg_15_53_inst : DFFX1 port map( D => n100, CLK => n4941, Q => 
                           RAM_15_53_port, QN => n_3023);
   RAM_reg_15_52_inst : DFFX1 port map( D => n99, CLK => n4941, Q => 
                           RAM_15_52_port, QN => n_3024);
   RAM_reg_15_51_inst : DFFX1 port map( D => n98, CLK => n4941, Q => 
                           RAM_15_51_port, QN => n_3025);
   RAM_reg_15_50_inst : DFFX1 port map( D => n97, CLK => n4941, Q => 
                           RAM_15_50_port, QN => n_3026);
   RAM_reg_15_49_inst : DFFX1 port map( D => n96, CLK => n4941, Q => 
                           RAM_15_49_port, QN => n_3027);
   RAM_reg_15_48_inst : DFFX1 port map( D => n95, CLK => n4941, Q => 
                           RAM_15_48_port, QN => n_3028);
   RAM_reg_15_47_inst : DFFX1 port map( D => n94, CLK => n4941, Q => 
                           RAM_15_47_port, QN => n_3029);
   RAM_reg_15_46_inst : DFFX1 port map( D => n93, CLK => n4941, Q => 
                           RAM_15_46_port, QN => n_3030);
   RAM_reg_15_45_inst : DFFX1 port map( D => n92, CLK => n4941, Q => 
                           RAM_15_45_port, QN => n_3031);
   RAM_reg_15_44_inst : DFFX1 port map( D => n91, CLK => n4941, Q => 
                           RAM_15_44_port, QN => n_3032);
   RAM_reg_15_43_inst : DFFX1 port map( D => n90, CLK => n4942, Q => 
                           RAM_15_43_port, QN => n_3033);
   RAM_reg_15_42_inst : DFFX1 port map( D => n89, CLK => n4942, Q => 
                           RAM_15_42_port, QN => n_3034);
   RAM_reg_15_41_inst : DFFX1 port map( D => n88, CLK => n4942, Q => 
                           RAM_15_41_port, QN => n_3035);
   RAM_reg_15_40_inst : DFFX1 port map( D => n87, CLK => n4942, Q => 
                           RAM_15_40_port, QN => n_3036);
   RAM_reg_15_39_inst : DFFX1 port map( D => n86, CLK => n4942, Q => 
                           RAM_15_39_port, QN => n_3037);
   RAM_reg_15_38_inst : DFFX1 port map( D => n85, CLK => n4942, Q => 
                           RAM_15_38_port, QN => n_3038);
   RAM_reg_15_37_inst : DFFX1 port map( D => n84, CLK => n4942, Q => 
                           RAM_15_37_port, QN => n_3039);
   RAM_reg_15_36_inst : DFFX1 port map( D => n83, CLK => n4942, Q => 
                           RAM_15_36_port, QN => n_3040);
   RAM_reg_15_35_inst : DFFX1 port map( D => n82, CLK => n4936, Q => 
                           RAM_15_35_port, QN => n_3041);
   RAM_reg_15_34_inst : DFFX1 port map( D => n81, CLK => n4936, Q => 
                           RAM_15_34_port, QN => n_3042);
   RAM_reg_15_33_inst : DFFX1 port map( D => n80, CLK => n4936, Q => 
                           RAM_15_33_port, QN => n_3043);
   RAM_reg_15_32_inst : DFFX1 port map( D => n79, CLK => n4936, Q => 
                           RAM_15_32_port, QN => n_3044);
   RAM_reg_15_31_inst : DFFX1 port map( D => n78, CLK => n4937, Q => 
                           RAM_15_31_port, QN => n_3045);
   RAM_reg_15_30_inst : DFFX1 port map( D => n77, CLK => n4937, Q => 
                           RAM_15_30_port, QN => n_3046);
   RAM_reg_15_29_inst : DFFX1 port map( D => n76, CLK => n4937, Q => 
                           RAM_15_29_port, QN => n_3047);
   RAM_reg_15_28_inst : DFFX1 port map( D => n75, CLK => n4937, Q => 
                           RAM_15_28_port, QN => n_3048);
   RAM_reg_15_27_inst : DFFX1 port map( D => n74, CLK => n4937, Q => 
                           RAM_15_27_port, QN => n_3049);
   RAM_reg_15_26_inst : DFFX1 port map( D => n73, CLK => n4937, Q => 
                           RAM_15_26_port, QN => n_3050);
   RAM_reg_15_25_inst : DFFX1 port map( D => n72, CLK => n4937, Q => 
                           RAM_15_25_port, QN => n_3051);
   RAM_reg_15_24_inst : DFFX1 port map( D => n71, CLK => n4937, Q => 
                           RAM_15_24_port, QN => n_3052);
   RAM_reg_15_23_inst : DFFX1 port map( D => n70, CLK => n4937, Q => 
                           RAM_15_23_port, QN => n_3053);
   RAM_reg_15_22_inst : DFFX1 port map( D => n69, CLK => n4937, Q => 
                           RAM_15_22_port, QN => n_3054);
   RAM_reg_15_21_inst : DFFX1 port map( D => n68, CLK => n4937, Q => 
                           RAM_15_21_port, QN => n_3055);
   RAM_reg_15_20_inst : DFFX1 port map( D => n67, CLK => n4937, Q => 
                           RAM_15_20_port, QN => n_3056);
   RAM_reg_15_19_inst : DFFX1 port map( D => n66, CLK => n4938, Q => 
                           RAM_15_19_port, QN => n_3057);
   RAM_reg_15_18_inst : DFFX1 port map( D => n65, CLK => n4938, Q => 
                           RAM_15_18_port, QN => n_3058);
   RAM_reg_15_17_inst : DFFX1 port map( D => n64, CLK => n4938, Q => 
                           RAM_15_17_port, QN => n_3059);
   RAM_reg_15_16_inst : DFFX1 port map( D => n63, CLK => n4938, Q => 
                           RAM_15_16_port, QN => n_3060);
   RAM_reg_15_15_inst : DFFX1 port map( D => n62, CLK => n4938, Q => 
                           RAM_15_15_port, QN => n_3061);
   RAM_reg_15_14_inst : DFFX1 port map( D => n61, CLK => n4938, Q => 
                           RAM_15_14_port, QN => n_3062);
   RAM_reg_15_13_inst : DFFX1 port map( D => n60, CLK => n4938, Q => 
                           RAM_15_13_port, QN => n_3063);
   RAM_reg_15_12_inst : DFFX1 port map( D => n59, CLK => n4938, Q => 
                           RAM_15_12_port, QN => n_3064);
   RAM_reg_15_11_inst : DFFX1 port map( D => n58, CLK => n4938, Q => 
                           RAM_15_11_port, QN => n_3065);
   RAM_reg_15_10_inst : DFFX1 port map( D => n57, CLK => n4938, Q => 
                           RAM_15_10_port, QN => n_3066);
   RAM_reg_15_9_inst : DFFX1 port map( D => n56, CLK => n4938, Q => 
                           RAM_15_9_port, QN => n_3067);
   RAM_reg_15_8_inst : DFFX1 port map( D => n55, CLK => n4938, Q => 
                           RAM_15_8_port, QN => n_3068);
   RAM_reg_15_7_inst : DFFX1 port map( D => n54, CLK => n4939, Q => 
                           RAM_15_7_port, QN => n_3069);
   RAM_reg_15_6_inst : DFFX1 port map( D => n53, CLK => n4939, Q => 
                           RAM_15_6_port, QN => n_3070);
   RAM_reg_15_5_inst : DFFX1 port map( D => n52, CLK => n4939, Q => 
                           RAM_15_5_port, QN => n_3071);
   RAM_reg_15_4_inst : DFFX1 port map( D => n51, CLK => n4939, Q => 
                           RAM_15_4_port, QN => n_3072);
   RAM_reg_15_3_inst : DFFX1 port map( D => n50, CLK => n4939, Q => 
                           RAM_15_3_port, QN => n_3073);
   RAM_reg_15_2_inst : DFFX1 port map( D => n49, CLK => n4939, Q => 
                           RAM_15_2_port, QN => n_3074);
   RAM_reg_15_1_inst : DFFX1 port map( D => n48, CLK => n4939, Q => 
                           RAM_15_1_port, QN => n_3075);
   RAM_reg_15_0_inst : DFFX1 port map( D => n47, CLK => n4939, Q => 
                           RAM_15_0_port, QN => n_3076);
   U43 : AO22X1 port map( IN1 => RAMDIN1(0), IN2 => n5608, IN3 => RAM_15_0_port
                           , IN4 => n5589, Q => n47);
   U44 : AO22X1 port map( IN1 => n5591, IN2 => RAMDIN1(1), IN3 => RAM_15_1_port
                           , IN4 => n5589, Q => n48);
   U45 : AO22X1 port map( IN1 => RAMDIN1(2), IN2 => n5590, IN3 => RAM_15_2_port
                           , IN4 => n5589, Q => n49);
   U46 : AO22X1 port map( IN1 => RAMDIN1(3), IN2 => n5591, IN3 => RAM_15_3_port
                           , IN4 => n5589, Q => n50);
   U47 : AO22X1 port map( IN1 => n5614, IN2 => RAMDIN1(4), IN3 => RAM_15_4_port
                           , IN4 => n5589, Q => n51);
   U48 : AO22X1 port map( IN1 => n5612, IN2 => RAMDIN1(5), IN3 => RAM_15_5_port
                           , IN4 => n5589, Q => n52);
   U49 : AO22X1 port map( IN1 => n5613, IN2 => RAMDIN1(6), IN3 => RAM_15_6_port
                           , IN4 => n5589, Q => n53);
   U50 : AO22X1 port map( IN1 => RAMDIN1(7), IN2 => n5614, IN3 => RAM_15_7_port
                           , IN4 => n5589, Q => n54);
   U51 : AO22X1 port map( IN1 => RAMDIN1(8), IN2 => n5612, IN3 => RAM_15_8_port
                           , IN4 => n5588, Q => n55);
   U52 : AO22X1 port map( IN1 => RAMDIN1(9), IN2 => n5612, IN3 => RAM_15_9_port
                           , IN4 => n5588, Q => n56);
   U53 : AO22X1 port map( IN1 => RAMDIN1(10), IN2 => n5614, IN3 => 
                           RAM_15_10_port, IN4 => n5588, Q => n57);
   U54 : AO22X1 port map( IN1 => RAMDIN1(11), IN2 => n5613, IN3 => 
                           RAM_15_11_port, IN4 => n5588, Q => n58);
   U55 : AO22X1 port map( IN1 => RAMDIN1(12), IN2 => n5613, IN3 => 
                           RAM_15_12_port, IN4 => n5588, Q => n59);
   U56 : AO22X1 port map( IN1 => RAMDIN1(13), IN2 => n5614, IN3 => 
                           RAM_15_13_port, IN4 => n5588, Q => n60);
   U57 : AO22X1 port map( IN1 => RAMDIN1(14), IN2 => n5592, IN3 => 
                           RAM_15_14_port, IN4 => n5588, Q => n61);
   U58 : AO22X1 port map( IN1 => RAMDIN1(15), IN2 => n5592, IN3 => 
                           RAM_15_15_port, IN4 => n5588, Q => n62);
   U59 : AO22X1 port map( IN1 => RAMDIN1(16), IN2 => n5592, IN3 => 
                           RAM_15_16_port, IN4 => n5588, Q => n63);
   U60 : AO22X1 port map( IN1 => RAMDIN1(17), IN2 => n5592, IN3 => 
                           RAM_15_17_port, IN4 => n5588, Q => n64);
   U61 : AO22X1 port map( IN1 => RAMDIN1(18), IN2 => n5592, IN3 => 
                           RAM_15_18_port, IN4 => n5588, Q => n65);
   U62 : AO22X1 port map( IN1 => n5593, IN2 => RAMDIN1(19), IN3 => 
                           RAM_15_19_port, IN4 => n5588, Q => n66);
   U63 : AO22X1 port map( IN1 => RAMDIN1(20), IN2 => n5593, IN3 => 
                           RAM_15_20_port, IN4 => n5587, Q => n67);
   U64 : AO22X1 port map( IN1 => RAMDIN1(21), IN2 => n5593, IN3 => 
                           RAM_15_21_port, IN4 => n5587, Q => n68);
   U65 : AO22X1 port map( IN1 => n2248, IN2 => n5593, IN3 => RAM_15_22_port, 
                           IN4 => n5587, Q => n69);
   U66 : AO22X1 port map( IN1 => RAMDIN1(23), IN2 => n5593, IN3 => 
                           RAM_15_23_port, IN4 => n5587, Q => n70);
   U67 : AO22X1 port map( IN1 => n2200, IN2 => n5594, IN3 => RAM_15_24_port, 
                           IN4 => n5587, Q => n71);
   U68 : AO22X1 port map( IN1 => RAMDIN1(25), IN2 => n5594, IN3 => 
                           RAM_15_25_port, IN4 => n5587, Q => n72);
   U69 : AO22X1 port map( IN1 => RAMDIN1(26), IN2 => n5594, IN3 => 
                           RAM_15_26_port, IN4 => n5587, Q => n73);
   U70 : AO22X1 port map( IN1 => RAMDIN1(27), IN2 => n5594, IN3 => 
                           RAM_15_27_port, IN4 => n5587, Q => n74);
   U71 : AO22X1 port map( IN1 => RAMDIN1(28), IN2 => n5594, IN3 => 
                           RAM_15_28_port, IN4 => n5587, Q => n75);
   U72 : AO22X1 port map( IN1 => RAMDIN1(29), IN2 => n5595, IN3 => 
                           RAM_15_29_port, IN4 => n5587, Q => n76);
   U73 : AO22X1 port map( IN1 => RAMDIN1(30), IN2 => n5595, IN3 => 
                           RAM_15_30_port, IN4 => n5587, Q => n77);
   U74 : AO22X1 port map( IN1 => n5595, IN2 => RAMDIN1(31), IN3 => 
                           RAM_15_31_port, IN4 => n5587, Q => n78);
   U75 : AO22X1 port map( IN1 => RAMDIN1(32), IN2 => n5595, IN3 => 
                           RAM_15_32_port, IN4 => n5586, Q => n79);
   U76 : AO22X1 port map( IN1 => RAMDIN1(33), IN2 => n5595, IN3 => 
                           RAM_15_33_port, IN4 => n5586, Q => n80);
   U77 : AO22X1 port map( IN1 => RAMDIN1(34), IN2 => n5596, IN3 => 
                           RAM_15_34_port, IN4 => n5586, Q => n81);
   U78 : AO22X1 port map( IN1 => n5596, IN2 => RAMDIN1(35), IN3 => 
                           RAM_15_35_port, IN4 => n5586, Q => n82);
   U79 : AO22X1 port map( IN1 => n5596, IN2 => RAMDIN1(36), IN3 => 
                           RAM_15_36_port, IN4 => n5586, Q => n83);
   U80 : AO22X1 port map( IN1 => n2558, IN2 => n5596, IN3 => RAM_15_37_port, 
                           IN4 => n5586, Q => n84);
   U81 : AO22X1 port map( IN1 => RAMDIN1(38), IN2 => n5596, IN3 => 
                           RAM_15_38_port, IN4 => n5586, Q => n85);
   U82 : AO22X1 port map( IN1 => n5597, IN2 => RAMDIN1(39), IN3 => 
                           RAM_15_39_port, IN4 => n5586, Q => n86);
   U83 : AO22X1 port map( IN1 => RAMDIN1(40), IN2 => n5597, IN3 => 
                           RAM_15_40_port, IN4 => n5586, Q => n87);
   U84 : AO22X1 port map( IN1 => n2507, IN2 => n5597, IN3 => RAM_15_41_port, 
                           IN4 => n5586, Q => n88);
   U85 : AO22X1 port map( IN1 => RAMDIN1(42), IN2 => n5597, IN3 => 
                           RAM_15_42_port, IN4 => n5586, Q => n89);
   U86 : AO22X1 port map( IN1 => n2560, IN2 => n5597, IN3 => RAM_15_43_port, 
                           IN4 => n5586, Q => n90);
   U87 : AO22X1 port map( IN1 => RAMDIN1(44), IN2 => n5598, IN3 => 
                           RAM_15_44_port, IN4 => n5585, Q => n91);
   U88 : AO22X1 port map( IN1 => RAMDIN1(45), IN2 => n5598, IN3 => 
                           RAM_15_45_port, IN4 => n5585, Q => n92);
   U89 : AO22X1 port map( IN1 => RAMDIN1(46), IN2 => n5598, IN3 => 
                           RAM_15_46_port, IN4 => n5585, Q => n93);
   U90 : AO22X1 port map( IN1 => RAMDIN1(47), IN2 => n5598, IN3 => 
                           RAM_15_47_port, IN4 => n5585, Q => n94);
   U91 : AO22X1 port map( IN1 => n2127, IN2 => n5598, IN3 => RAM_15_48_port, 
                           IN4 => n5585, Q => n95);
   U92 : AO22X1 port map( IN1 => RAMDIN1(49), IN2 => n5599, IN3 => 
                           RAM_15_49_port, IN4 => n5585, Q => n96);
   U93 : AO22X1 port map( IN1 => RAMDIN1(50), IN2 => n5599, IN3 => 
                           RAM_15_50_port, IN4 => n5585, Q => n97);
   U94 : AO22X1 port map( IN1 => RAMDIN1(51), IN2 => n5599, IN3 => 
                           RAM_15_51_port, IN4 => n5585, Q => n98);
   U95 : AO22X1 port map( IN1 => n2555, IN2 => n5599, IN3 => RAM_15_52_port, 
                           IN4 => n5585, Q => n99);
   U96 : AO22X1 port map( IN1 => n5599, IN2 => RAMDIN1(53), IN3 => 
                           RAM_15_53_port, IN4 => n5585, Q => n100);
   U97 : AO22X1 port map( IN1 => RAMDIN1(54), IN2 => n5600, IN3 => 
                           RAM_15_54_port, IN4 => n5585, Q => n101);
   U98 : AO22X1 port map( IN1 => RAMDIN1(55), IN2 => n5600, IN3 => 
                           RAM_15_55_port, IN4 => n5585, Q => n102);
   U102 : AO22X1 port map( IN1 => RAMDIN1(59), IN2 => n5601, IN3 => 
                           RAM_15_59_port, IN4 => n5584, Q => n106);
   U103 : AO22X1 port map( IN1 => RAMDIN1(60), IN2 => n5601, IN3 => 
                           RAM_15_60_port, IN4 => n5584, Q => n107);
   U104 : AO22X1 port map( IN1 => RAMDIN1(61), IN2 => n5601, IN3 => 
                           RAM_15_61_port, IN4 => n5584, Q => n108);
   U105 : AO22X1 port map( IN1 => RAMDIN1(62), IN2 => n5601, IN3 => 
                           RAM_15_62_port, IN4 => n5584, Q => n109);
   U106 : AO22X1 port map( IN1 => RAMDIN1(63), IN2 => n5601, IN3 => 
                           RAM_15_63_port, IN4 => n5584, Q => n110);
   U107 : AO22X1 port map( IN1 => n5602, IN2 => RAMDIN1(64), IN3 => 
                           RAM_15_64_port, IN4 => n5584, Q => n111);
   U108 : AO22X1 port map( IN1 => RAMDIN1(65), IN2 => n5602, IN3 => 
                           RAM_15_65_port, IN4 => n5584, Q => n112);
   U109 : AO22X1 port map( IN1 => RAMDIN1(66), IN2 => n5602, IN3 => 
                           RAM_15_66_port, IN4 => n5584, Q => n113);
   U110 : AO22X1 port map( IN1 => RAMDIN1(67), IN2 => n5602, IN3 => 
                           RAM_15_67_port, IN4 => n5584, Q => n114);
   U111 : AO22X1 port map( IN1 => RAMDIN1(68), IN2 => n5602, IN3 => 
                           RAM_15_68_port, IN4 => n5583, Q => n115);
   U112 : AO22X1 port map( IN1 => n5603, IN2 => RAMDIN1(69), IN3 => 
                           RAM_15_69_port, IN4 => n5583, Q => n116);
   U113 : AO22X1 port map( IN1 => n5603, IN2 => RAMDIN1(70), IN3 => 
                           RAM_15_70_port, IN4 => n5583, Q => n117);
   U114 : AO22X1 port map( IN1 => n5603, IN2 => RAMDIN1(71), IN3 => 
                           RAM_15_71_port, IN4 => n5583, Q => n118);
   U115 : AO22X1 port map( IN1 => RAMDIN1(72), IN2 => n5603, IN3 => 
                           RAM_15_72_port, IN4 => n5583, Q => n119);
   U116 : AO22X1 port map( IN1 => RAMDIN1(73), IN2 => n5603, IN3 => 
                           RAM_15_73_port, IN4 => n5583, Q => n120);
   U117 : AO22X1 port map( IN1 => RAMDIN1(74), IN2 => n5604, IN3 => 
                           RAM_15_74_port, IN4 => n5583, Q => n121);
   U118 : AO22X1 port map( IN1 => RAMDIN1(75), IN2 => n5604, IN3 => 
                           RAM_15_75_port, IN4 => n5583, Q => n122);
   U119 : AO22X1 port map( IN1 => RAMDIN1(76), IN2 => n5604, IN3 => 
                           RAM_15_76_port, IN4 => n5583, Q => n123);
   U120 : AO22X1 port map( IN1 => RAMDIN1(77), IN2 => n5604, IN3 => 
                           RAM_15_77_port, IN4 => n5583, Q => n124);
   U121 : AO22X1 port map( IN1 => RAMDIN1(78), IN2 => n5604, IN3 => 
                           RAM_15_78_port, IN4 => n5583, Q => n125);
   U122 : AO22X1 port map( IN1 => RAMDIN1(79), IN2 => n5605, IN3 => 
                           RAM_15_79_port, IN4 => n5583, Q => n126);
   U123 : AO22X1 port map( IN1 => RAMDIN1(80), IN2 => n5605, IN3 => 
                           RAM_15_80_port, IN4 => n5582, Q => n127);
   U124 : AO22X1 port map( IN1 => RAMDIN1(81), IN2 => n5605, IN3 => 
                           RAM_15_81_port, IN4 => n5582, Q => n128);
   U125 : AO22X1 port map( IN1 => RAMDIN1(82), IN2 => n5605, IN3 => 
                           RAM_15_82_port, IN4 => n5582, Q => n129);
   U126 : AO22X1 port map( IN1 => RAMDIN1(83), IN2 => n5605, IN3 => 
                           RAM_15_83_port, IN4 => n5582, Q => n130);
   U127 : AO22X1 port map( IN1 => RAMDIN1(84), IN2 => n5606, IN3 => 
                           RAM_15_84_port, IN4 => n5582, Q => n131);
   U128 : AO22X1 port map( IN1 => RAMDIN1(85), IN2 => n5606, IN3 => 
                           RAM_15_85_port, IN4 => n5582, Q => n132);
   U129 : AO22X1 port map( IN1 => RAMDIN1(86), IN2 => n5606, IN3 => 
                           RAM_15_86_port, IN4 => n5582, Q => n133);
   U130 : AO22X1 port map( IN1 => RAMDIN1(87), IN2 => n5606, IN3 => 
                           RAM_15_87_port, IN4 => n5582, Q => n134);
   U131 : AO22X1 port map( IN1 => RAMDIN1(88), IN2 => n5606, IN3 => 
                           RAM_15_88_port, IN4 => n5582, Q => n135);
   U132 : AO22X1 port map( IN1 => RAMDIN1(89), IN2 => n5607, IN3 => 
                           RAM_15_89_port, IN4 => n5582, Q => n136);
   U133 : AO22X1 port map( IN1 => RAMDIN1(90), IN2 => n5607, IN3 => 
                           RAM_15_90_port, IN4 => n5582, Q => n137);
   U134 : AO22X1 port map( IN1 => RAMDIN1(91), IN2 => n5607, IN3 => 
                           RAM_15_91_port, IN4 => n5582, Q => n138);
   U135 : AO22X1 port map( IN1 => RAMDIN1(92), IN2 => n5607, IN3 => 
                           RAM_15_92_port, IN4 => n5581, Q => n139);
   U136 : AO22X1 port map( IN1 => RAMDIN1(93), IN2 => n5607, IN3 => 
                           RAM_15_93_port, IN4 => n5581, Q => n140);
   U137 : AO22X1 port map( IN1 => RAMDIN1(94), IN2 => n5608, IN3 => 
                           RAM_15_94_port, IN4 => n5581, Q => n141);
   U138 : AO22X1 port map( IN1 => RAMDIN1(95), IN2 => n5608, IN3 => 
                           RAM_15_95_port, IN4 => n5581, Q => n142);
   U139 : AO22X1 port map( IN1 => n5608, IN2 => RAMDIN1(96), IN3 => 
                           RAM_15_96_port, IN4 => n5581, Q => n143);
   U140 : AO22X1 port map( IN1 => n5608, IN2 => RAMDIN1(97), IN3 => 
                           RAM_15_97_port, IN4 => n5581, Q => n144);
   U141 : AO22X1 port map( IN1 => n5608, IN2 => RAMDIN1(98), IN3 => 
                           RAM_15_98_port, IN4 => n5581, Q => n145);
   U142 : AO22X1 port map( IN1 => n2503, IN2 => n5609, IN3 => RAM_15_99_port, 
                           IN4 => n5581, Q => n146);
   U143 : AO22X1 port map( IN1 => n5609, IN2 => RAMDIN1(100), IN3 => 
                           RAM_15_100_port, IN4 => n5581, Q => n147);
   U144 : AO22X1 port map( IN1 => n5609, IN2 => RAMDIN1(101), IN3 => 
                           RAM_15_101_port, IN4 => n5581, Q => n148);
   U145 : AO22X1 port map( IN1 => n5609, IN2 => RAMDIN1(102), IN3 => 
                           RAM_15_102_port, IN4 => n5581, Q => n149);
   U146 : AO22X1 port map( IN1 => RAMDIN1(103), IN2 => n5609, IN3 => 
                           RAM_15_103_port, IN4 => n5581, Q => n150);
   U147 : AO22X1 port map( IN1 => n5610, IN2 => RAMDIN1(104), IN3 => 
                           RAM_15_104_port, IN4 => n5580, Q => n151);
   U148 : AO22X1 port map( IN1 => n5610, IN2 => RAMDIN1(105), IN3 => 
                           RAM_15_105_port, IN4 => n5580, Q => n152);
   U149 : AO22X1 port map( IN1 => RAMDIN1(106), IN2 => n5610, IN3 => 
                           RAM_15_106_port, IN4 => n5580, Q => n153);
   U150 : AO22X1 port map( IN1 => RAMDIN1(107), IN2 => n5610, IN3 => 
                           RAM_15_107_port, IN4 => n5580, Q => n154);
   U151 : AO22X1 port map( IN1 => RAMDIN1(108), IN2 => n5610, IN3 => 
                           RAM_15_108_port, IN4 => n5580, Q => n155);
   U152 : AO22X1 port map( IN1 => RAMDIN1(109), IN2 => n5611, IN3 => 
                           RAM_15_109_port, IN4 => n5580, Q => n156);
   U153 : AO22X1 port map( IN1 => RAMDIN1(110), IN2 => n5611, IN3 => 
                           RAM_15_110_port, IN4 => n5580, Q => n157);
   U154 : AO22X1 port map( IN1 => RAMDIN1(111), IN2 => n5611, IN3 => 
                           RAM_15_111_port, IN4 => n5580, Q => n158);
   U155 : AO22X1 port map( IN1 => RAMDIN1(112), IN2 => n5611, IN3 => 
                           RAM_15_112_port, IN4 => n5580, Q => n159);
   U156 : AO22X1 port map( IN1 => RAMDIN1(113), IN2 => n5611, IN3 => 
                           RAM_15_113_port, IN4 => n5580, Q => n160);
   U157 : AO22X1 port map( IN1 => RAMDIN1(114), IN2 => n5612, IN3 => 
                           RAM_15_114_port, IN4 => n5580, Q => n161);
   U158 : AO22X1 port map( IN1 => RAMDIN1(115), IN2 => n5612, IN3 => 
                           RAM_15_115_port, IN4 => n5580, Q => n162);
   U159 : AO22X1 port map( IN1 => RAMDIN1(116), IN2 => n5612, IN3 => 
                           RAM_15_116_port, IN4 => n5579, Q => n163);
   U160 : AO22X1 port map( IN1 => n5612, IN2 => RAMDIN1(117), IN3 => 
                           RAM_15_117_port, IN4 => n5579, Q => n164);
   U161 : AO22X1 port map( IN1 => n5612, IN2 => RAMDIN1(118), IN3 => 
                           RAM_15_118_port, IN4 => n5579, Q => n165);
   U162 : AO22X1 port map( IN1 => n5613, IN2 => RAMDIN1(119), IN3 => 
                           RAM_15_119_port, IN4 => n5579, Q => n166);
   U163 : AO22X1 port map( IN1 => RAMDIN1(120), IN2 => n5613, IN3 => 
                           RAM_15_120_port, IN4 => n5579, Q => n167);
   U164 : AO22X1 port map( IN1 => RAMDIN1(121), IN2 => n5613, IN3 => 
                           RAM_15_121_port, IN4 => n5579, Q => n168);
   U165 : AO22X1 port map( IN1 => RAMDIN1(122), IN2 => n5613, IN3 => 
                           RAM_15_122_port, IN4 => n5579, Q => n169);
   U166 : AO22X1 port map( IN1 => RAMDIN1(123), IN2 => n5613, IN3 => 
                           RAM_15_123_port, IN4 => n5579, Q => n170);
   U167 : AO22X1 port map( IN1 => RAMDIN1(124), IN2 => n5614, IN3 => 
                           RAM_15_124_port, IN4 => n5579, Q => n171);
   U168 : AO22X1 port map( IN1 => RAMDIN1(125), IN2 => n5614, IN3 => 
                           RAM_15_125_port, IN4 => n5579, Q => n172);
   U169 : AO22X1 port map( IN1 => RAMDIN1(126), IN2 => n5614, IN3 => 
                           RAM_15_126_port, IN4 => n5579, Q => n173);
   U170 : AO22X1 port map( IN1 => RAMDIN1(127), IN2 => n5614, IN3 => 
                           RAM_15_127_port, IN4 => n5579, Q => n174);
   U171 : AO22X1 port map( IN1 => n5558, IN2 => RAMDIN1(0), IN3 => 
                           RAM_14_0_port, IN4 => n5547, Q => n175);
   U172 : AO22X1 port map( IN1 => n5559, IN2 => RAMDIN1(1), IN3 => 
                           RAM_14_1_port, IN4 => n5547, Q => n176);
   U173 : AO22X1 port map( IN1 => n5548, IN2 => RAMDIN1(2), IN3 => 
                           RAM_14_2_port, IN4 => n5547, Q => n177);
   U174 : AO22X1 port map( IN1 => n5548, IN2 => RAMDIN1(3), IN3 => 
                           RAM_14_3_port, IN4 => n5547, Q => n178);
   U175 : AO22X1 port map( IN1 => n5570, IN2 => RAMDIN1(4), IN3 => 
                           RAM_14_4_port, IN4 => n5547, Q => n179);
   U176 : AO22X1 port map( IN1 => n5572, IN2 => RAMDIN1(5), IN3 => 
                           RAM_14_5_port, IN4 => n5547, Q => n180);
   U177 : AO22X1 port map( IN1 => n5571, IN2 => RAMDIN1(6), IN3 => 
                           RAM_14_6_port, IN4 => n5547, Q => n181);
   U178 : AO22X1 port map( IN1 => n5570, IN2 => RAMDIN1(7), IN3 => 
                           RAM_14_7_port, IN4 => n5547, Q => n182);
   U179 : AO22X1 port map( IN1 => n5572, IN2 => RAMDIN1(8), IN3 => 
                           RAM_14_8_port, IN4 => n5546, Q => n183);
   U180 : AO22X1 port map( IN1 => n5572, IN2 => RAMDIN1(9), IN3 => 
                           RAM_14_9_port, IN4 => n5546, Q => n184);
   U181 : AO22X1 port map( IN1 => n5571, IN2 => RAMDIN1(10), IN3 => 
                           RAM_14_10_port, IN4 => n5546, Q => n185);
   U182 : AO22X1 port map( IN1 => n5570, IN2 => RAMDIN1(11), IN3 => 
                           RAM_14_11_port, IN4 => n5546, Q => n186);
   U183 : AO22X1 port map( IN1 => n5572, IN2 => RAMDIN1(12), IN3 => 
                           RAM_14_12_port, IN4 => n5546, Q => n187);
   U184 : AO22X1 port map( IN1 => RAMDIN1(13), IN2 => n5571, IN3 => 
                           RAM_14_13_port, IN4 => n5546, Q => n188);
   U185 : AO22X1 port map( IN1 => RAMDIN1(14), IN2 => n5550, IN3 => 
                           RAM_14_14_port, IN4 => n5546, Q => n189);
   U186 : AO22X1 port map( IN1 => n5550, IN2 => RAMDIN1(15), IN3 => 
                           RAM_14_15_port, IN4 => n5546, Q => n190);
   U187 : AO22X1 port map( IN1 => RAMDIN1(16), IN2 => n5550, IN3 => 
                           RAM_14_16_port, IN4 => n5546, Q => n191);
   U188 : AO22X1 port map( IN1 => n5550, IN2 => RAMDIN1(17), IN3 => 
                           RAM_14_17_port, IN4 => n5546, Q => n192);
   U189 : AO22X1 port map( IN1 => n5550, IN2 => RAMDIN1(18), IN3 => 
                           RAM_14_18_port, IN4 => n5546, Q => n193);
   U190 : AO22X1 port map( IN1 => n5551, IN2 => RAMDIN1(19), IN3 => 
                           RAM_14_19_port, IN4 => n5546, Q => n194);
   U191 : AO22X1 port map( IN1 => n5551, IN2 => RAMDIN1(20), IN3 => 
                           RAM_14_20_port, IN4 => n5545, Q => n195);
   U192 : AO22X1 port map( IN1 => n5551, IN2 => RAMDIN1(21), IN3 => 
                           RAM_14_21_port, IN4 => n5545, Q => n196);
   U193 : AO22X1 port map( IN1 => n5551, IN2 => n2248, IN3 => RAM_14_22_port, 
                           IN4 => n5545, Q => n197);
   U194 : AO22X1 port map( IN1 => n5551, IN2 => RAMDIN1(23), IN3 => 
                           RAM_14_23_port, IN4 => n5545, Q => n198);
   U195 : AO22X1 port map( IN1 => n5552, IN2 => n2201, IN3 => RAM_14_24_port, 
                           IN4 => n5545, Q => n199);
   U196 : AO22X1 port map( IN1 => n5552, IN2 => RAMDIN1(25), IN3 => 
                           RAM_14_25_port, IN4 => n5545, Q => n200);
   U197 : AO22X1 port map( IN1 => n5552, IN2 => RAMDIN1(26), IN3 => 
                           RAM_14_26_port, IN4 => n5545, Q => n201);
   U198 : AO22X1 port map( IN1 => n5552, IN2 => RAMDIN1(27), IN3 => 
                           RAM_14_27_port, IN4 => n5545, Q => n202);
   U199 : AO22X1 port map( IN1 => RAMDIN1(28), IN2 => n5552, IN3 => 
                           RAM_14_28_port, IN4 => n5545, Q => n203);
   U200 : AO22X1 port map( IN1 => n5553, IN2 => RAMDIN1(29), IN3 => 
                           RAM_14_29_port, IN4 => n5545, Q => n204);
   U201 : AO22X1 port map( IN1 => n5553, IN2 => RAMDIN1(30), IN3 => 
                           RAM_14_30_port, IN4 => n5545, Q => n205);
   U202 : AO22X1 port map( IN1 => n5553, IN2 => RAMDIN1(31), IN3 => 
                           RAM_14_31_port, IN4 => n5545, Q => n206);
   U203 : AO22X1 port map( IN1 => n5553, IN2 => RAMDIN1(32), IN3 => 
                           RAM_14_32_port, IN4 => n5544, Q => n207);
   U204 : AO22X1 port map( IN1 => n5553, IN2 => RAMDIN1(33), IN3 => 
                           RAM_14_33_port, IN4 => n5544, Q => n208);
   U205 : AO22X1 port map( IN1 => n5554, IN2 => RAMDIN1(34), IN3 => 
                           RAM_14_34_port, IN4 => n5544, Q => n209);
   U206 : AO22X1 port map( IN1 => n5554, IN2 => RAMDIN1(35), IN3 => 
                           RAM_14_35_port, IN4 => n5544, Q => n210);
   U207 : AO22X1 port map( IN1 => n5554, IN2 => RAMDIN1(36), IN3 => 
                           RAM_14_36_port, IN4 => n5544, Q => n211);
   U208 : AO22X1 port map( IN1 => n5554, IN2 => n2559, IN3 => RAM_14_37_port, 
                           IN4 => n5544, Q => n212);
   U209 : AO22X1 port map( IN1 => n5554, IN2 => RAMDIN1(38), IN3 => 
                           RAM_14_38_port, IN4 => n5544, Q => n213);
   U210 : AO22X1 port map( IN1 => n5555, IN2 => RAMDIN1(39), IN3 => 
                           RAM_14_39_port, IN4 => n5544, Q => n214);
   U211 : AO22X1 port map( IN1 => n5555, IN2 => RAMDIN1(40), IN3 => 
                           RAM_14_40_port, IN4 => n5544, Q => n215);
   U212 : AO22X1 port map( IN1 => n5555, IN2 => n2506, IN3 => RAM_14_41_port, 
                           IN4 => n5544, Q => n216);
   U213 : AO22X1 port map( IN1 => n5555, IN2 => RAMDIN1(42), IN3 => 
                           RAM_14_42_port, IN4 => n5544, Q => n217);
   U214 : AO22X1 port map( IN1 => n5555, IN2 => n2560, IN3 => RAM_14_43_port, 
                           IN4 => n5544, Q => n218);
   U215 : AO22X1 port map( IN1 => n5556, IN2 => RAMDIN1(44), IN3 => 
                           RAM_14_44_port, IN4 => n5543, Q => n219);
   U216 : AO22X1 port map( IN1 => n5556, IN2 => RAMDIN1(45), IN3 => 
                           RAM_14_45_port, IN4 => n5543, Q => n220);
   U217 : AO22X1 port map( IN1 => RAMDIN1(46), IN2 => n5556, IN3 => 
                           RAM_14_46_port, IN4 => n5543, Q => n221);
   U218 : AO22X1 port map( IN1 => n5556, IN2 => RAMDIN1(47), IN3 => 
                           RAM_14_47_port, IN4 => n5543, Q => n222);
   U219 : AO22X1 port map( IN1 => n5556, IN2 => n2127, IN3 => RAM_14_48_port, 
                           IN4 => n5543, Q => n223);
   U220 : AO22X1 port map( IN1 => n5557, IN2 => RAMDIN1(49), IN3 => 
                           RAM_14_49_port, IN4 => n5543, Q => n224);
   U221 : AO22X1 port map( IN1 => n5557, IN2 => RAMDIN1(50), IN3 => 
                           RAM_14_50_port, IN4 => n5543, Q => n225);
   U222 : AO22X1 port map( IN1 => n5557, IN2 => RAMDIN1(51), IN3 => 
                           RAM_14_51_port, IN4 => n5543, Q => n226);
   U223 : AO22X1 port map( IN1 => n5557, IN2 => n2, IN3 => RAM_14_52_port, IN4 
                           => n5543, Q => n227);
   U224 : AO22X1 port map( IN1 => n5557, IN2 => RAMDIN1(53), IN3 => 
                           RAM_14_53_port, IN4 => n5543, Q => n228);
   U225 : AO22X1 port map( IN1 => n5558, IN2 => RAMDIN1(54), IN3 => 
                           RAM_14_54_port, IN4 => n5543, Q => n229);
   U226 : AO22X1 port map( IN1 => n5558, IN2 => RAMDIN1(55), IN3 => 
                           RAM_14_55_port, IN4 => n5543, Q => n230);
   U239 : AO22X1 port map( IN1 => n5560, IN2 => RAMDIN1(68), IN3 => 
                           RAM_14_68_port, IN4 => n5541, Q => n243);
   U240 : AO22X1 port map( IN1 => n5561, IN2 => RAMDIN1(69), IN3 => 
                           RAM_14_69_port, IN4 => n5541, Q => n244);
   U241 : AO22X1 port map( IN1 => n5561, IN2 => RAMDIN1(70), IN3 => 
                           RAM_14_70_port, IN4 => n5541, Q => n245);
   U242 : AO22X1 port map( IN1 => n5561, IN2 => RAMDIN1(71), IN3 => 
                           RAM_14_71_port, IN4 => n5541, Q => n246);
   U243 : AO22X1 port map( IN1 => n5561, IN2 => RAMDIN1(72), IN3 => 
                           RAM_14_72_port, IN4 => n5541, Q => n247);
   U244 : AO22X1 port map( IN1 => RAMDIN1(73), IN2 => n5561, IN3 => 
                           RAM_14_73_port, IN4 => n5541, Q => n248);
   U245 : AO22X1 port map( IN1 => n5562, IN2 => RAMDIN1(74), IN3 => 
                           RAM_14_74_port, IN4 => n5541, Q => n249);
   U246 : AO22X1 port map( IN1 => n5562, IN2 => RAMDIN1(75), IN3 => 
                           RAM_14_75_port, IN4 => n5541, Q => n250);
   U247 : AO22X1 port map( IN1 => n5562, IN2 => RAMDIN1(76), IN3 => 
                           RAM_14_76_port, IN4 => n5541, Q => n251);
   U248 : AO22X1 port map( IN1 => n5562, IN2 => RAMDIN1(77), IN3 => 
                           RAM_14_77_port, IN4 => n5541, Q => n252);
   U249 : AO22X1 port map( IN1 => n5562, IN2 => RAMDIN1(78), IN3 => 
                           RAM_14_78_port, IN4 => n5541, Q => n253);
   U250 : AO22X1 port map( IN1 => RAMDIN1(79), IN2 => n5563, IN3 => 
                           RAM_14_79_port, IN4 => n5541, Q => n254);
   U251 : AO22X1 port map( IN1 => RAMDIN1(80), IN2 => n5563, IN3 => 
                           RAM_14_80_port, IN4 => n5540, Q => n255);
   U252 : AO22X1 port map( IN1 => n5563, IN2 => RAMDIN1(81), IN3 => 
                           RAM_14_81_port, IN4 => n5540, Q => n256);
   U253 : AO22X1 port map( IN1 => n5563, IN2 => RAMDIN1(82), IN3 => 
                           RAM_14_82_port, IN4 => n5540, Q => n257);
   U254 : AO22X1 port map( IN1 => n5563, IN2 => RAMDIN1(83), IN3 => 
                           RAM_14_83_port, IN4 => n5540, Q => n258);
   U255 : AO22X1 port map( IN1 => n5564, IN2 => RAMDIN1(84), IN3 => 
                           RAM_14_84_port, IN4 => n5540, Q => n259);
   U256 : AO22X1 port map( IN1 => n5564, IN2 => RAMDIN1(85), IN3 => 
                           RAM_14_85_port, IN4 => n5540, Q => n260);
   U257 : AO22X1 port map( IN1 => n5564, IN2 => RAMDIN1(86), IN3 => 
                           RAM_14_86_port, IN4 => n5540, Q => n261);
   U258 : AO22X1 port map( IN1 => n5564, IN2 => RAMDIN1(87), IN3 => 
                           RAM_14_87_port, IN4 => n5540, Q => n262);
   U259 : AO22X1 port map( IN1 => RAMDIN1(88), IN2 => n5564, IN3 => 
                           RAM_14_88_port, IN4 => n5540, Q => n263);
   U260 : AO22X1 port map( IN1 => n5565, IN2 => RAMDIN1(89), IN3 => 
                           RAM_14_89_port, IN4 => n5540, Q => n264);
   U261 : AO22X1 port map( IN1 => n5565, IN2 => RAMDIN1(90), IN3 => 
                           RAM_14_90_port, IN4 => n5540, Q => n265);
   U262 : AO22X1 port map( IN1 => n5565, IN2 => RAMDIN1(91), IN3 => 
                           RAM_14_91_port, IN4 => n5540, Q => n266);
   U263 : AO22X1 port map( IN1 => n5565, IN2 => RAMDIN1(92), IN3 => 
                           RAM_14_92_port, IN4 => n5539, Q => n267);
   U264 : AO22X1 port map( IN1 => n5565, IN2 => RAMDIN1(93), IN3 => 
                           RAM_14_93_port, IN4 => n5539, Q => n268);
   U265 : AO22X1 port map( IN1 => n5566, IN2 => RAMDIN1(94), IN3 => 
                           RAM_14_94_port, IN4 => n5539, Q => n269);
   U266 : AO22X1 port map( IN1 => n5566, IN2 => RAMDIN1(95), IN3 => 
                           RAM_14_95_port, IN4 => n5539, Q => n270);
   U267 : AO22X1 port map( IN1 => n5566, IN2 => RAMDIN1(96), IN3 => 
                           RAM_14_96_port, IN4 => n5539, Q => n271);
   U268 : AO22X1 port map( IN1 => n5566, IN2 => RAMDIN1(97), IN3 => 
                           RAM_14_97_port, IN4 => n5539, Q => n272);
   U269 : AO22X1 port map( IN1 => n5566, IN2 => RAMDIN1(98), IN3 => 
                           RAM_14_98_port, IN4 => n5539, Q => n273);
   U270 : AO22X1 port map( IN1 => n5567, IN2 => n2502, IN3 => RAM_14_99_port, 
                           IN4 => n5539, Q => n274);
   U271 : AO22X1 port map( IN1 => n5567, IN2 => RAMDIN1(100), IN3 => 
                           RAM_14_100_port, IN4 => n5539, Q => n275);
   U272 : AO22X1 port map( IN1 => n5567, IN2 => RAMDIN1(101), IN3 => 
                           RAM_14_101_port, IN4 => n5539, Q => n276);
   U273 : AO22X1 port map( IN1 => n5567, IN2 => RAMDIN1(102), IN3 => 
                           RAM_14_102_port, IN4 => n5539, Q => n277);
   U274 : AO22X1 port map( IN1 => n5567, IN2 => RAMDIN1(103), IN3 => 
                           RAM_14_103_port, IN4 => n5539, Q => n278);
   U275 : AO22X1 port map( IN1 => n5568, IN2 => RAMDIN1(104), IN3 => 
                           RAM_14_104_port, IN4 => n5538, Q => n279);
   U276 : AO22X1 port map( IN1 => n5568, IN2 => RAMDIN1(105), IN3 => 
                           RAM_14_105_port, IN4 => n5538, Q => n280);
   U277 : AO22X1 port map( IN1 => n5568, IN2 => RAMDIN1(106), IN3 => 
                           RAM_14_106_port, IN4 => n5538, Q => n281);
   U278 : AO22X1 port map( IN1 => n5568, IN2 => RAMDIN1(107), IN3 => 
                           RAM_14_107_port, IN4 => n5538, Q => n282);
   U279 : AO22X1 port map( IN1 => n5568, IN2 => RAMDIN1(108), IN3 => 
                           RAM_14_108_port, IN4 => n5538, Q => n283);
   U280 : AO22X1 port map( IN1 => n5569, IN2 => RAMDIN1(109), IN3 => 
                           RAM_14_109_port, IN4 => n5538, Q => n284);
   U281 : AO22X1 port map( IN1 => RAMDIN1(110), IN2 => n5569, IN3 => 
                           RAM_14_110_port, IN4 => n5538, Q => n285);
   U282 : AO22X1 port map( IN1 => n5569, IN2 => RAMDIN1(111), IN3 => 
                           RAM_14_111_port, IN4 => n5538, Q => n286);
   U283 : AO22X1 port map( IN1 => RAMDIN1(112), IN2 => n5569, IN3 => 
                           RAM_14_112_port, IN4 => n5538, Q => n287);
   U284 : AO22X1 port map( IN1 => n5569, IN2 => RAMDIN1(113), IN3 => 
                           RAM_14_113_port, IN4 => n5538, Q => n288);
   U285 : AO22X1 port map( IN1 => n5570, IN2 => RAMDIN1(114), IN3 => 
                           RAM_14_114_port, IN4 => n5538, Q => n289);
   U286 : AO22X1 port map( IN1 => n5570, IN2 => RAMDIN1(115), IN3 => 
                           RAM_14_115_port, IN4 => n5538, Q => n290);
   U287 : AO22X1 port map( IN1 => n5570, IN2 => RAMDIN1(116), IN3 => 
                           RAM_14_116_port, IN4 => n5537, Q => n291);
   U288 : AO22X1 port map( IN1 => n5570, IN2 => RAMDIN1(117), IN3 => 
                           RAM_14_117_port, IN4 => n5537, Q => n292);
   U289 : AO22X1 port map( IN1 => n5570, IN2 => RAMDIN1(118), IN3 => 
                           RAM_14_118_port, IN4 => n5537, Q => n293);
   U290 : AO22X1 port map( IN1 => n5571, IN2 => RAMDIN1(119), IN3 => 
                           RAM_14_119_port, IN4 => n5537, Q => n294);
   U291 : AO22X1 port map( IN1 => n5571, IN2 => RAMDIN1(120), IN3 => 
                           RAM_14_120_port, IN4 => n5537, Q => n295);
   U292 : AO22X1 port map( IN1 => n5571, IN2 => RAMDIN1(121), IN3 => 
                           RAM_14_121_port, IN4 => n5537, Q => n296);
   U293 : AO22X1 port map( IN1 => n5571, IN2 => RAMDIN1(122), IN3 => 
                           RAM_14_122_port, IN4 => n5537, Q => n297);
   U294 : AO22X1 port map( IN1 => n5571, IN2 => RAMDIN1(123), IN3 => 
                           RAM_14_123_port, IN4 => n5537, Q => n298);
   U295 : AO22X1 port map( IN1 => n5572, IN2 => RAMDIN1(124), IN3 => 
                           RAM_14_124_port, IN4 => n5537, Q => n299);
   U296 : AO22X1 port map( IN1 => n5572, IN2 => RAMDIN1(125), IN3 => 
                           RAM_14_125_port, IN4 => n5537, Q => n300);
   U297 : AO22X1 port map( IN1 => n5572, IN2 => RAMDIN1(126), IN3 => 
                           RAM_14_126_port, IN4 => n5537, Q => n301);
   U298 : AO22X1 port map( IN1 => RAMDIN1(127), IN2 => n5572, IN3 => 
                           RAM_14_127_port, IN4 => n5537, Q => n302);
   U299 : AO22X1 port map( IN1 => n5509, IN2 => RAMDIN1(0), IN3 => 
                           RAM_13_0_port, IN4 => n5505, Q => n303);
   U300 : AO22X1 port map( IN1 => n5508, IN2 => RAMDIN1(1), IN3 => 
                           RAM_13_1_port, IN4 => n5505, Q => n304);
   U301 : AO22X1 port map( IN1 => n5506, IN2 => RAMDIN1(2), IN3 => 
                           RAM_13_2_port, IN4 => n5505, Q => n305);
   U302 : AO22X1 port map( IN1 => n5506, IN2 => RAMDIN1(3), IN3 => 
                           RAM_13_3_port, IN4 => n5505, Q => n306);
   U303 : AO22X1 port map( IN1 => n5528, IN2 => RAMDIN1(4), IN3 => 
                           RAM_13_4_port, IN4 => n5505, Q => n307);
   U304 : AO22X1 port map( IN1 => n5528, IN2 => RAMDIN1(5), IN3 => 
                           RAM_13_5_port, IN4 => n5505, Q => n308);
   U305 : AO22X1 port map( IN1 => n5529, IN2 => RAMDIN1(6), IN3 => 
                           RAM_13_6_port, IN4 => n5505, Q => n309);
   U306 : AO22X1 port map( IN1 => n5530, IN2 => RAMDIN1(7), IN3 => 
                           RAM_13_7_port, IN4 => n5505, Q => n310);
   U307 : AO22X1 port map( IN1 => n5530, IN2 => RAMDIN1(8), IN3 => 
                           RAM_13_8_port, IN4 => n5504, Q => n311);
   U308 : AO22X1 port map( IN1 => n5530, IN2 => RAMDIN1(9), IN3 => 
                           RAM_13_9_port, IN4 => n5504, Q => n312);
   U309 : AO22X1 port map( IN1 => n5529, IN2 => RAMDIN1(10), IN3 => 
                           RAM_13_10_port, IN4 => n5504, Q => n313);
   U310 : AO22X1 port map( IN1 => n5528, IN2 => RAMDIN1(11), IN3 => 
                           RAM_13_11_port, IN4 => n5504, Q => n314);
   U311 : AO22X1 port map( IN1 => n5530, IN2 => RAMDIN1(12), IN3 => 
                           RAM_13_12_port, IN4 => n5504, Q => n315);
   U312 : AO22X1 port map( IN1 => RAMDIN1(13), IN2 => n5529, IN3 => 
                           RAM_13_13_port, IN4 => n5504, Q => n316);
   U313 : AO22X1 port map( IN1 => RAMDIN1(14), IN2 => n5508, IN3 => 
                           RAM_13_14_port, IN4 => n5504, Q => n317);
   U314 : AO22X1 port map( IN1 => n5508, IN2 => RAMDIN1(15), IN3 => 
                           RAM_13_15_port, IN4 => n5504, Q => n318);
   U315 : AO22X1 port map( IN1 => RAMDIN1(16), IN2 => n5508, IN3 => 
                           RAM_13_16_port, IN4 => n5504, Q => n319);
   U316 : AO22X1 port map( IN1 => n5508, IN2 => RAMDIN1(17), IN3 => 
                           RAM_13_17_port, IN4 => n5504, Q => n320);
   U317 : AO22X1 port map( IN1 => n5508, IN2 => RAMDIN1(18), IN3 => 
                           RAM_13_18_port, IN4 => n5504, Q => n321);
   U318 : AO22X1 port map( IN1 => n5509, IN2 => RAMDIN1(19), IN3 => 
                           RAM_13_19_port, IN4 => n5504, Q => n322);
   U319 : AO22X1 port map( IN1 => n5509, IN2 => RAMDIN1(20), IN3 => 
                           RAM_13_20_port, IN4 => n5503, Q => n323);
   U320 : AO22X1 port map( IN1 => RAMDIN1(21), IN2 => n5509, IN3 => 
                           RAM_13_21_port, IN4 => n5503, Q => n324);
   U321 : AO22X1 port map( IN1 => n5509, IN2 => n2248, IN3 => RAM_13_22_port, 
                           IN4 => n5503, Q => n325);
   U322 : AO22X1 port map( IN1 => n5509, IN2 => RAMDIN1(23), IN3 => 
                           RAM_13_23_port, IN4 => n5503, Q => n326);
   U323 : AO22X1 port map( IN1 => n5510, IN2 => n2201, IN3 => RAM_13_24_port, 
                           IN4 => n5503, Q => n327);
   U324 : AO22X1 port map( IN1 => n5510, IN2 => RAMDIN1(25), IN3 => 
                           RAM_13_25_port, IN4 => n5503, Q => n328);
   U325 : AO22X1 port map( IN1 => n5510, IN2 => RAMDIN1(26), IN3 => 
                           RAM_13_26_port, IN4 => n5503, Q => n329);
   U326 : AO22X1 port map( IN1 => n5510, IN2 => RAMDIN1(27), IN3 => 
                           RAM_13_27_port, IN4 => n5503, Q => n330);
   U327 : AO22X1 port map( IN1 => RAMDIN1(28), IN2 => n5510, IN3 => 
                           RAM_13_28_port, IN4 => n5503, Q => n331);
   U328 : AO22X1 port map( IN1 => n5511, IN2 => RAMDIN1(29), IN3 => 
                           RAM_13_29_port, IN4 => n5503, Q => n332);
   U329 : AO22X1 port map( IN1 => n5511, IN2 => RAMDIN1(30), IN3 => 
                           RAM_13_30_port, IN4 => n5503, Q => n333);
   U330 : AO22X1 port map( IN1 => n5511, IN2 => RAMDIN1(31), IN3 => 
                           RAM_13_31_port, IN4 => n5503, Q => n334);
   U331 : AO22X1 port map( IN1 => n5511, IN2 => RAMDIN1(32), IN3 => 
                           RAM_13_32_port, IN4 => n5502, Q => n335);
   U332 : AO22X1 port map( IN1 => n5511, IN2 => RAMDIN1(33), IN3 => 
                           RAM_13_33_port, IN4 => n5502, Q => n336);
   U333 : AO22X1 port map( IN1 => n5512, IN2 => RAMDIN1(34), IN3 => 
                           RAM_13_34_port, IN4 => n5502, Q => n337);
   U334 : AO22X1 port map( IN1 => n5512, IN2 => RAMDIN1(35), IN3 => 
                           RAM_13_35_port, IN4 => n5502, Q => n338);
   U335 : AO22X1 port map( IN1 => n5512, IN2 => RAMDIN1(36), IN3 => 
                           RAM_13_36_port, IN4 => n5502, Q => n339);
   U336 : AO22X1 port map( IN1 => n5512, IN2 => n2559, IN3 => RAM_13_37_port, 
                           IN4 => n5502, Q => n340);
   U337 : AO22X1 port map( IN1 => n5512, IN2 => RAMDIN1(38), IN3 => 
                           RAM_13_38_port, IN4 => n5502, Q => n341);
   U338 : AO22X1 port map( IN1 => n5513, IN2 => RAMDIN1(39), IN3 => 
                           RAM_13_39_port, IN4 => n5502, Q => n342);
   U339 : AO22X1 port map( IN1 => n5513, IN2 => RAMDIN1(40), IN3 => 
                           RAM_13_40_port, IN4 => n5502, Q => n343);
   U340 : AO22X1 port map( IN1 => n5513, IN2 => n2507, IN3 => RAM_13_41_port, 
                           IN4 => n5502, Q => n344);
   U341 : AO22X1 port map( IN1 => n5513, IN2 => RAMDIN1(42), IN3 => 
                           RAM_13_42_port, IN4 => n5502, Q => n345);
   U342 : AO22X1 port map( IN1 => n5513, IN2 => n2560, IN3 => RAM_13_43_port, 
                           IN4 => n5502, Q => n346);
   U343 : AO22X1 port map( IN1 => RAMDIN1(44), IN2 => n5514, IN3 => 
                           RAM_13_44_port, IN4 => n5501, Q => n347);
   U344 : AO22X1 port map( IN1 => RAMDIN1(45), IN2 => n5514, IN3 => 
                           RAM_13_45_port, IN4 => n5501, Q => n348);
   U345 : AO22X1 port map( IN1 => RAMDIN1(46), IN2 => n5514, IN3 => 
                           RAM_13_46_port, IN4 => n5501, Q => n349);
   U346 : AO22X1 port map( IN1 => n5514, IN2 => RAMDIN1(47), IN3 => 
                           RAM_13_47_port, IN4 => n5501, Q => n350);
   U347 : AO22X1 port map( IN1 => n5514, IN2 => n2127, IN3 => RAM_13_48_port, 
                           IN4 => n5501, Q => n351);
   U348 : AO22X1 port map( IN1 => n5515, IN2 => RAMDIN1(49), IN3 => 
                           RAM_13_49_port, IN4 => n5501, Q => n352);
   U349 : AO22X1 port map( IN1 => n5515, IN2 => RAMDIN1(50), IN3 => 
                           RAM_13_50_port, IN4 => n5501, Q => n353);
   U350 : AO22X1 port map( IN1 => n5515, IN2 => RAMDIN1(51), IN3 => 
                           RAM_13_51_port, IN4 => n5501, Q => n354);
   U351 : AO22X1 port map( IN1 => n5515, IN2 => n2555, IN3 => RAM_13_52_port, 
                           IN4 => n5501, Q => n355);
   U352 : AO22X1 port map( IN1 => n5515, IN2 => RAMDIN1(53), IN3 => 
                           RAM_13_53_port, IN4 => n5501, Q => n356);
   U353 : AO22X1 port map( IN1 => n5516, IN2 => RAMDIN1(54), IN3 => 
                           RAM_13_54_port, IN4 => n5501, Q => n357);
   U354 : AO22X1 port map( IN1 => n5516, IN2 => RAMDIN1(55), IN3 => 
                           RAM_13_55_port, IN4 => n5501, Q => n358);
   U355 : AO22X1 port map( IN1 => n5516, IN2 => RAMDIN1(56), IN3 => 
                           RAM_13_56_port, IN4 => n5500, Q => n359);
   U356 : AO22X1 port map( IN1 => n5516, IN2 => RAMDIN1(57), IN3 => 
                           RAM_13_57_port, IN4 => n5500, Q => n360);
   U357 : AO22X1 port map( IN1 => n5516, IN2 => RAMDIN1(58), IN3 => 
                           RAM_13_58_port, IN4 => n5500, Q => n361);
   U358 : AO22X1 port map( IN1 => n5517, IN2 => RAMDIN1(59), IN3 => 
                           RAM_13_59_port, IN4 => n5500, Q => n362);
   U359 : AO22X1 port map( IN1 => n5517, IN2 => RAMDIN1(60), IN3 => 
                           RAM_13_60_port, IN4 => n5500, Q => n363);
   U360 : AO22X1 port map( IN1 => n5517, IN2 => RAMDIN1(61), IN3 => 
                           RAM_13_61_port, IN4 => n5500, Q => n364);
   U361 : AO22X1 port map( IN1 => n5517, IN2 => RAMDIN1(62), IN3 => 
                           RAM_13_62_port, IN4 => n5500, Q => n365);
   U362 : AO22X1 port map( IN1 => n5517, IN2 => RAMDIN1(63), IN3 => 
                           RAM_13_63_port, IN4 => n5500, Q => n366);
   U363 : AO22X1 port map( IN1 => n5518, IN2 => RAMDIN1(64), IN3 => 
                           RAM_13_64_port, IN4 => n5500, Q => n367);
   U364 : AO22X1 port map( IN1 => n5518, IN2 => RAMDIN1(65), IN3 => 
                           RAM_13_65_port, IN4 => n5500, Q => n368);
   U365 : AO22X1 port map( IN1 => n5518, IN2 => RAMDIN1(66), IN3 => 
                           RAM_13_66_port, IN4 => n5500, Q => n369);
   U366 : AO22X1 port map( IN1 => n5518, IN2 => RAMDIN1(67), IN3 => 
                           RAM_13_67_port, IN4 => n5500, Q => n370);
   U367 : AO22X1 port map( IN1 => n5518, IN2 => RAMDIN1(68), IN3 => 
                           RAM_13_68_port, IN4 => n5499, Q => n371);
   U368 : AO22X1 port map( IN1 => RAMDIN1(69), IN2 => n5519, IN3 => 
                           RAM_13_69_port, IN4 => n5499, Q => n372);
   U369 : AO22X1 port map( IN1 => n5519, IN2 => RAMDIN1(70), IN3 => 
                           RAM_13_70_port, IN4 => n5499, Q => n373);
   U370 : AO22X1 port map( IN1 => n5519, IN2 => RAMDIN1(71), IN3 => 
                           RAM_13_71_port, IN4 => n5499, Q => n374);
   U371 : AO22X1 port map( IN1 => n5519, IN2 => RAMDIN1(72), IN3 => 
                           RAM_13_72_port, IN4 => n5499, Q => n375);
   U372 : AO22X1 port map( IN1 => n5519, IN2 => RAMDIN1(73), IN3 => 
                           RAM_13_73_port, IN4 => n5499, Q => n376);
   U373 : AO22X1 port map( IN1 => n5520, IN2 => RAMDIN1(74), IN3 => 
                           RAM_13_74_port, IN4 => n5499, Q => n377);
   U374 : AO22X1 port map( IN1 => n5520, IN2 => RAMDIN1(75), IN3 => 
                           RAM_13_75_port, IN4 => n5499, Q => n378);
   U375 : AO22X1 port map( IN1 => n5520, IN2 => RAMDIN1(76), IN3 => 
                           RAM_13_76_port, IN4 => n5499, Q => n379);
   U376 : AO22X1 port map( IN1 => n5520, IN2 => RAMDIN1(77), IN3 => 
                           RAM_13_77_port, IN4 => n5499, Q => n380);
   U377 : AO22X1 port map( IN1 => n5520, IN2 => RAMDIN1(78), IN3 => 
                           RAM_13_78_port, IN4 => n5499, Q => n381);
   U378 : AO22X1 port map( IN1 => n5521, IN2 => RAMDIN1(79), IN3 => 
                           RAM_13_79_port, IN4 => n5499, Q => n382);
   U379 : AO22X1 port map( IN1 => RAMDIN1(80), IN2 => n5521, IN3 => 
                           RAM_13_80_port, IN4 => n5498, Q => n383);
   U380 : AO22X1 port map( IN1 => n5521, IN2 => RAMDIN1(81), IN3 => 
                           RAM_13_81_port, IN4 => n5498, Q => n384);
   U381 : AO22X1 port map( IN1 => n5521, IN2 => RAMDIN1(82), IN3 => 
                           RAM_13_82_port, IN4 => n5498, Q => n385);
   U382 : AO22X1 port map( IN1 => n5521, IN2 => RAMDIN1(83), IN3 => 
                           RAM_13_83_port, IN4 => n5498, Q => n386);
   U383 : AO22X1 port map( IN1 => n5522, IN2 => RAMDIN1(84), IN3 => 
                           RAM_13_84_port, IN4 => n5498, Q => n387);
   U384 : AO22X1 port map( IN1 => n5522, IN2 => RAMDIN1(85), IN3 => 
                           RAM_13_85_port, IN4 => n5498, Q => n388);
   U385 : AO22X1 port map( IN1 => n5522, IN2 => RAMDIN1(86), IN3 => 
                           RAM_13_86_port, IN4 => n5498, Q => n389);
   U386 : AO22X1 port map( IN1 => n5522, IN2 => RAMDIN1(87), IN3 => 
                           RAM_13_87_port, IN4 => n5498, Q => n390);
   U387 : AO22X1 port map( IN1 => RAMDIN1(88), IN2 => n5522, IN3 => 
                           RAM_13_88_port, IN4 => n5498, Q => n391);
   U388 : AO22X1 port map( IN1 => n5523, IN2 => RAMDIN1(89), IN3 => 
                           RAM_13_89_port, IN4 => n5498, Q => n392);
   U389 : AO22X1 port map( IN1 => n5523, IN2 => RAMDIN1(90), IN3 => 
                           RAM_13_90_port, IN4 => n5498, Q => n393);
   U390 : AO22X1 port map( IN1 => n5523, IN2 => RAMDIN1(91), IN3 => 
                           RAM_13_91_port, IN4 => n5498, Q => n394);
   U391 : AO22X1 port map( IN1 => n5523, IN2 => RAMDIN1(92), IN3 => 
                           RAM_13_92_port, IN4 => n5497, Q => n395);
   U392 : AO22X1 port map( IN1 => n5523, IN2 => RAMDIN1(93), IN3 => 
                           RAM_13_93_port, IN4 => n5497, Q => n396);
   U393 : AO22X1 port map( IN1 => n5524, IN2 => RAMDIN1(94), IN3 => 
                           RAM_13_94_port, IN4 => n5497, Q => n397);
   U394 : AO22X1 port map( IN1 => n5524, IN2 => RAMDIN1(95), IN3 => 
                           RAM_13_95_port, IN4 => n5497, Q => n398);
   U395 : AO22X1 port map( IN1 => n5524, IN2 => RAMDIN1(96), IN3 => 
                           RAM_13_96_port, IN4 => n5497, Q => n399);
   U396 : AO22X1 port map( IN1 => RAMDIN1(97), IN2 => n5524, IN3 => 
                           RAM_13_97_port, IN4 => n5497, Q => n400);
   U397 : AO22X1 port map( IN1 => n5524, IN2 => RAMDIN1(98), IN3 => 
                           RAM_13_98_port, IN4 => n5497, Q => n401);
   U398 : AO22X1 port map( IN1 => n5525, IN2 => n2503, IN3 => RAM_13_99_port, 
                           IN4 => n5497, Q => n402);
   U399 : AO22X1 port map( IN1 => n5525, IN2 => RAMDIN1(100), IN3 => 
                           RAM_13_100_port, IN4 => n5497, Q => n403);
   U400 : AO22X1 port map( IN1 => n5525, IN2 => RAMDIN1(101), IN3 => 
                           RAM_13_101_port, IN4 => n5497, Q => n404);
   U401 : AO22X1 port map( IN1 => n5525, IN2 => RAMDIN1(102), IN3 => 
                           RAM_13_102_port, IN4 => n5497, Q => n405);
   U402 : AO22X1 port map( IN1 => n5525, IN2 => RAMDIN1(103), IN3 => 
                           RAM_13_103_port, IN4 => n5497, Q => n406);
   U403 : AO22X1 port map( IN1 => n5526, IN2 => RAMDIN1(104), IN3 => 
                           RAM_13_104_port, IN4 => n5496, Q => n407);
   U404 : AO22X1 port map( IN1 => n5526, IN2 => RAMDIN1(105), IN3 => 
                           RAM_13_105_port, IN4 => n5496, Q => n408);
   U405 : AO22X1 port map( IN1 => n5526, IN2 => RAMDIN1(106), IN3 => 
                           RAM_13_106_port, IN4 => n5496, Q => n409);
   U406 : AO22X1 port map( IN1 => n5526, IN2 => RAMDIN1(107), IN3 => 
                           RAM_13_107_port, IN4 => n5496, Q => n410);
   U407 : AO22X1 port map( IN1 => n5526, IN2 => RAMDIN1(108), IN3 => 
                           RAM_13_108_port, IN4 => n5496, Q => n411);
   U408 : AO22X1 port map( IN1 => n5527, IN2 => RAMDIN1(109), IN3 => 
                           RAM_13_109_port, IN4 => n5496, Q => n412);
   U409 : AO22X1 port map( IN1 => RAMDIN1(110), IN2 => n5527, IN3 => 
                           RAM_13_110_port, IN4 => n5496, Q => n413);
   U410 : AO22X1 port map( IN1 => n5527, IN2 => RAMDIN1(111), IN3 => 
                           RAM_13_111_port, IN4 => n5496, Q => n414);
   U411 : AO22X1 port map( IN1 => RAMDIN1(112), IN2 => n5527, IN3 => 
                           RAM_13_112_port, IN4 => n5496, Q => n415);
   U412 : AO22X1 port map( IN1 => n5527, IN2 => RAMDIN1(113), IN3 => 
                           RAM_13_113_port, IN4 => n5496, Q => n416);
   U413 : AO22X1 port map( IN1 => n5528, IN2 => RAMDIN1(114), IN3 => 
                           RAM_13_114_port, IN4 => n5496, Q => n417);
   U414 : AO22X1 port map( IN1 => n5528, IN2 => RAMDIN1(115), IN3 => 
                           RAM_13_115_port, IN4 => n5496, Q => n418);
   U415 : AO22X1 port map( IN1 => n5528, IN2 => RAMDIN1(116), IN3 => 
                           RAM_13_116_port, IN4 => n5495, Q => n419);
   U416 : AO22X1 port map( IN1 => n5528, IN2 => RAMDIN1(117), IN3 => 
                           RAM_13_117_port, IN4 => n5495, Q => n420);
   U417 : AO22X1 port map( IN1 => n5528, IN2 => RAMDIN1(118), IN3 => 
                           RAM_13_118_port, IN4 => n5495, Q => n421);
   U418 : AO22X1 port map( IN1 => n5529, IN2 => RAMDIN1(119), IN3 => 
                           RAM_13_119_port, IN4 => n5495, Q => n422);
   U419 : AO22X1 port map( IN1 => n5529, IN2 => RAMDIN1(120), IN3 => 
                           RAM_13_120_port, IN4 => n5495, Q => n423);
   U420 : AO22X1 port map( IN1 => n5529, IN2 => RAMDIN1(121), IN3 => 
                           RAM_13_121_port, IN4 => n5495, Q => n424);
   U421 : AO22X1 port map( IN1 => n5529, IN2 => RAMDIN1(122), IN3 => 
                           RAM_13_122_port, IN4 => n5495, Q => n425);
   U422 : AO22X1 port map( IN1 => n5529, IN2 => RAMDIN1(123), IN3 => 
                           RAM_13_123_port, IN4 => n5495, Q => n426);
   U423 : AO22X1 port map( IN1 => n5530, IN2 => RAMDIN1(124), IN3 => 
                           RAM_13_124_port, IN4 => n5495, Q => n427);
   U424 : AO22X1 port map( IN1 => n5530, IN2 => RAMDIN1(125), IN3 => 
                           RAM_13_125_port, IN4 => n5495, Q => n428);
   U425 : AO22X1 port map( IN1 => n5530, IN2 => RAMDIN1(126), IN3 => 
                           RAM_13_126_port, IN4 => n5495, Q => n429);
   U426 : AO22X1 port map( IN1 => RAMDIN1(127), IN2 => n5530, IN3 => 
                           RAM_13_127_port, IN4 => n5495, Q => n430);
   U427 : AO22X1 port map( IN1 => n5467, IN2 => RAMDIN1(0), IN3 => 
                           RAM_12_0_port, IN4 => n5463, Q => n431);
   U428 : AO22X1 port map( IN1 => n5466, IN2 => RAMDIN1(1), IN3 => 
                           RAM_12_1_port, IN4 => n5463, Q => n432);
   U429 : AO22X1 port map( IN1 => n5464, IN2 => RAMDIN1(2), IN3 => 
                           RAM_12_2_port, IN4 => n5463, Q => n433);
   U430 : AO22X1 port map( IN1 => n5464, IN2 => RAMDIN1(3), IN3 => 
                           RAM_12_3_port, IN4 => n5463, Q => n434);
   U431 : AO22X1 port map( IN1 => n5486, IN2 => RAMDIN1(4), IN3 => 
                           RAM_12_4_port, IN4 => n5463, Q => n435);
   U432 : AO22X1 port map( IN1 => n5488, IN2 => RAMDIN1(5), IN3 => 
                           RAM_12_5_port, IN4 => n5463, Q => n436);
   U433 : AO22X1 port map( IN1 => n5487, IN2 => RAMDIN1(6), IN3 => 
                           RAM_12_6_port, IN4 => n5463, Q => n437);
   U434 : AO22X1 port map( IN1 => n5486, IN2 => RAMDIN1(7), IN3 => 
                           RAM_12_7_port, IN4 => n5463, Q => n438);
   U435 : AO22X1 port map( IN1 => RAMDIN1(8), IN2 => n5488, IN3 => 
                           RAM_12_8_port, IN4 => n5462, Q => n439);
   U436 : AO22X1 port map( IN1 => n5488, IN2 => RAMDIN1(9), IN3 => 
                           RAM_12_9_port, IN4 => n5462, Q => n440);
   U437 : AO22X1 port map( IN1 => n5487, IN2 => RAMDIN1(10), IN3 => 
                           RAM_12_10_port, IN4 => n5462, Q => n441);
   U438 : AO22X1 port map( IN1 => n5486, IN2 => RAMDIN1(11), IN3 => 
                           RAM_12_11_port, IN4 => n5462, Q => n442);
   U439 : AO22X1 port map( IN1 => n5488, IN2 => RAMDIN1(12), IN3 => 
                           RAM_12_12_port, IN4 => n5462, Q => n443);
   U440 : AO22X1 port map( IN1 => RAMDIN1(13), IN2 => n5487, IN3 => 
                           RAM_12_13_port, IN4 => n5462, Q => n444);
   U441 : AO22X1 port map( IN1 => RAMDIN1(14), IN2 => n5466, IN3 => 
                           RAM_12_14_port, IN4 => n5462, Q => n445);
   U442 : AO22X1 port map( IN1 => n5466, IN2 => RAMDIN1(15), IN3 => 
                           RAM_12_15_port, IN4 => n5462, Q => n446);
   U443 : AO22X1 port map( IN1 => RAMDIN1(16), IN2 => n5466, IN3 => 
                           RAM_12_16_port, IN4 => n5462, Q => n447);
   U444 : AO22X1 port map( IN1 => n5466, IN2 => RAMDIN1(17), IN3 => 
                           RAM_12_17_port, IN4 => n5462, Q => n448);
   U445 : AO22X1 port map( IN1 => n5466, IN2 => RAMDIN1(18), IN3 => 
                           RAM_12_18_port, IN4 => n5462, Q => n449);
   U446 : AO22X1 port map( IN1 => n5467, IN2 => RAMDIN1(19), IN3 => 
                           RAM_12_19_port, IN4 => n5462, Q => n450);
   U447 : AO22X1 port map( IN1 => n5467, IN2 => RAMDIN1(20), IN3 => 
                           RAM_12_20_port, IN4 => n5461, Q => n451);
   U448 : AO22X1 port map( IN1 => n5467, IN2 => RAMDIN1(21), IN3 => 
                           RAM_12_21_port, IN4 => n5461, Q => n452);
   U449 : AO22X1 port map( IN1 => n5467, IN2 => n2248, IN3 => RAM_12_22_port, 
                           IN4 => n5461, Q => n453);
   U450 : AO22X1 port map( IN1 => n5467, IN2 => RAMDIN1(23), IN3 => 
                           RAM_12_23_port, IN4 => n5461, Q => n454);
   U451 : AO22X1 port map( IN1 => n5468, IN2 => n2201, IN3 => RAM_12_24_port, 
                           IN4 => n5461, Q => n455);
   U452 : AO22X1 port map( IN1 => n5468, IN2 => RAMDIN1(25), IN3 => 
                           RAM_12_25_port, IN4 => n5461, Q => n456);
   U453 : AO22X1 port map( IN1 => n5468, IN2 => RAMDIN1(26), IN3 => 
                           RAM_12_26_port, IN4 => n5461, Q => n457);
   U454 : AO22X1 port map( IN1 => n5468, IN2 => RAMDIN1(27), IN3 => 
                           RAM_12_27_port, IN4 => n5461, Q => n458);
   U455 : AO22X1 port map( IN1 => RAMDIN1(28), IN2 => n5468, IN3 => 
                           RAM_12_28_port, IN4 => n5461, Q => n459);
   U456 : AO22X1 port map( IN1 => n5469, IN2 => RAMDIN1(29), IN3 => 
                           RAM_12_29_port, IN4 => n5461, Q => n460);
   U457 : AO22X1 port map( IN1 => n5469, IN2 => RAMDIN1(30), IN3 => 
                           RAM_12_30_port, IN4 => n5461, Q => n461);
   U458 : AO22X1 port map( IN1 => n5469, IN2 => RAMDIN1(31), IN3 => 
                           RAM_12_31_port, IN4 => n5461, Q => n462);
   U459 : AO22X1 port map( IN1 => n5469, IN2 => RAMDIN1(32), IN3 => 
                           RAM_12_32_port, IN4 => n5460, Q => n463);
   U460 : AO22X1 port map( IN1 => n5469, IN2 => RAMDIN1(33), IN3 => 
                           RAM_12_33_port, IN4 => n5460, Q => n464);
   U461 : AO22X1 port map( IN1 => n5470, IN2 => RAMDIN1(34), IN3 => 
                           RAM_12_34_port, IN4 => n5460, Q => n465);
   U462 : AO22X1 port map( IN1 => n5470, IN2 => RAMDIN1(35), IN3 => 
                           RAM_12_35_port, IN4 => n5460, Q => n466);
   U463 : AO22X1 port map( IN1 => n5470, IN2 => RAMDIN1(36), IN3 => 
                           RAM_12_36_port, IN4 => n5460, Q => n467);
   U464 : AO22X1 port map( IN1 => n5470, IN2 => n1, IN3 => RAM_12_37_port, IN4 
                           => n5460, Q => n468);
   U465 : AO22X1 port map( IN1 => n5470, IN2 => RAMDIN1(38), IN3 => 
                           RAM_12_38_port, IN4 => n5460, Q => n469);
   U466 : AO22X1 port map( IN1 => n5471, IN2 => RAMDIN1(39), IN3 => 
                           RAM_12_39_port, IN4 => n5460, Q => n470);
   U467 : AO22X1 port map( IN1 => n5471, IN2 => RAMDIN1(40), IN3 => 
                           RAM_12_40_port, IN4 => n5460, Q => n471);
   U468 : AO22X1 port map( IN1 => n5471, IN2 => n2507, IN3 => RAM_12_41_port, 
                           IN4 => n5460, Q => n472);
   U469 : AO22X1 port map( IN1 => n5471, IN2 => RAMDIN1(42), IN3 => 
                           RAM_12_42_port, IN4 => n5460, Q => n473);
   U470 : AO22X1 port map( IN1 => n5471, IN2 => n2561, IN3 => RAM_12_43_port, 
                           IN4 => n5460, Q => n474);
   U471 : AO22X1 port map( IN1 => RAMDIN1(44), IN2 => n5472, IN3 => 
                           RAM_12_44_port, IN4 => n5459, Q => n475);
   U472 : AO22X1 port map( IN1 => n5472, IN2 => RAMDIN1(45), IN3 => 
                           RAM_12_45_port, IN4 => n5459, Q => n476);
   U473 : AO22X1 port map( IN1 => RAMDIN1(46), IN2 => n5472, IN3 => 
                           RAM_12_46_port, IN4 => n5459, Q => n477);
   U474 : AO22X1 port map( IN1 => n5472, IN2 => RAMDIN1(47), IN3 => 
                           RAM_12_47_port, IN4 => n5459, Q => n478);
   U475 : AO22X1 port map( IN1 => n5472, IN2 => n2126, IN3 => RAM_12_48_port, 
                           IN4 => n5459, Q => n479);
   U476 : AO22X1 port map( IN1 => n5473, IN2 => RAMDIN1(49), IN3 => 
                           RAM_12_49_port, IN4 => n5459, Q => n480);
   U477 : AO22X1 port map( IN1 => n5473, IN2 => RAMDIN1(50), IN3 => 
                           RAM_12_50_port, IN4 => n5459, Q => n481);
   U478 : AO22X1 port map( IN1 => n5473, IN2 => RAMDIN1(51), IN3 => 
                           RAM_12_51_port, IN4 => n5459, Q => n482);
   U479 : AO22X1 port map( IN1 => n5473, IN2 => n2, IN3 => RAM_12_52_port, IN4 
                           => n5459, Q => n483);
   U480 : AO22X1 port map( IN1 => n5473, IN2 => RAMDIN1(53), IN3 => 
                           RAM_12_53_port, IN4 => n5459, Q => n484);
   U481 : AO22X1 port map( IN1 => n5474, IN2 => RAMDIN1(54), IN3 => 
                           RAM_12_54_port, IN4 => n5459, Q => n485);
   U482 : AO22X1 port map( IN1 => n5474, IN2 => RAMDIN1(55), IN3 => 
                           RAM_12_55_port, IN4 => n5459, Q => n486);
   U483 : AO22X1 port map( IN1 => n5474, IN2 => RAMDIN1(56), IN3 => 
                           RAM_12_56_port, IN4 => n5458, Q => n487);
   U484 : AO22X1 port map( IN1 => n5474, IN2 => RAMDIN1(57), IN3 => 
                           RAM_12_57_port, IN4 => n5458, Q => n488);
   U485 : AO22X1 port map( IN1 => n5474, IN2 => RAMDIN1(58), IN3 => 
                           RAM_12_58_port, IN4 => n5458, Q => n489);
   U486 : AO22X1 port map( IN1 => n5475, IN2 => RAMDIN1(59), IN3 => 
                           RAM_12_59_port, IN4 => n5458, Q => n490);
   U487 : AO22X1 port map( IN1 => n5475, IN2 => RAMDIN1(60), IN3 => 
                           RAM_12_60_port, IN4 => n5458, Q => n491);
   U488 : AO22X1 port map( IN1 => n5475, IN2 => RAMDIN1(61), IN3 => 
                           RAM_12_61_port, IN4 => n5458, Q => n492);
   U489 : AO22X1 port map( IN1 => n5475, IN2 => RAMDIN1(62), IN3 => 
                           RAM_12_62_port, IN4 => n5458, Q => n493);
   U490 : AO22X1 port map( IN1 => n5475, IN2 => RAMDIN1(63), IN3 => 
                           RAM_12_63_port, IN4 => n5458, Q => n494);
   U491 : AO22X1 port map( IN1 => n5476, IN2 => RAMDIN1(64), IN3 => 
                           RAM_12_64_port, IN4 => n5458, Q => n495);
   U492 : AO22X1 port map( IN1 => n5476, IN2 => RAMDIN1(65), IN3 => 
                           RAM_12_65_port, IN4 => n5458, Q => n496);
   U493 : AO22X1 port map( IN1 => n5476, IN2 => RAMDIN1(66), IN3 => 
                           RAM_12_66_port, IN4 => n5458, Q => n497);
   U494 : AO22X1 port map( IN1 => n5476, IN2 => RAMDIN1(67), IN3 => 
                           RAM_12_67_port, IN4 => n5458, Q => n498);
   U495 : AO22X1 port map( IN1 => n5476, IN2 => RAMDIN1(68), IN3 => 
                           RAM_12_68_port, IN4 => n5457, Q => n499);
   U496 : AO22X1 port map( IN1 => n5477, IN2 => RAMDIN1(69), IN3 => 
                           RAM_12_69_port, IN4 => n5457, Q => n500);
   U497 : AO22X1 port map( IN1 => n5477, IN2 => RAMDIN1(70), IN3 => 
                           RAM_12_70_port, IN4 => n5457, Q => n501);
   U498 : AO22X1 port map( IN1 => n5477, IN2 => RAMDIN1(71), IN3 => 
                           RAM_12_71_port, IN4 => n5457, Q => n502);
   U499 : AO22X1 port map( IN1 => n5477, IN2 => RAMDIN1(72), IN3 => 
                           RAM_12_72_port, IN4 => n5457, Q => n503);
   U500 : AO22X1 port map( IN1 => n5477, IN2 => RAMDIN1(73), IN3 => 
                           RAM_12_73_port, IN4 => n5457, Q => n504);
   U501 : AO22X1 port map( IN1 => n5478, IN2 => RAMDIN1(74), IN3 => 
                           RAM_12_74_port, IN4 => n5457, Q => n505);
   U502 : AO22X1 port map( IN1 => n5478, IN2 => RAMDIN1(75), IN3 => 
                           RAM_12_75_port, IN4 => n5457, Q => n506);
   U503 : AO22X1 port map( IN1 => n5478, IN2 => RAMDIN1(76), IN3 => 
                           RAM_12_76_port, IN4 => n5457, Q => n507);
   U504 : AO22X1 port map( IN1 => n5478, IN2 => RAMDIN1(77), IN3 => 
                           RAM_12_77_port, IN4 => n5457, Q => n508);
   U505 : AO22X1 port map( IN1 => n5478, IN2 => RAMDIN1(78), IN3 => 
                           RAM_12_78_port, IN4 => n5457, Q => n509);
   U506 : AO22X1 port map( IN1 => n5479, IN2 => RAMDIN1(79), IN3 => 
                           RAM_12_79_port, IN4 => n5457, Q => n510);
   U507 : AO22X1 port map( IN1 => RAMDIN1(80), IN2 => n5479, IN3 => 
                           RAM_12_80_port, IN4 => n5456, Q => n511);
   U508 : AO22X1 port map( IN1 => n5479, IN2 => RAMDIN1(81), IN3 => 
                           RAM_12_81_port, IN4 => n5456, Q => n512);
   U509 : AO22X1 port map( IN1 => n5479, IN2 => RAMDIN1(82), IN3 => 
                           RAM_12_82_port, IN4 => n5456, Q => n513);
   U510 : AO22X1 port map( IN1 => n5479, IN2 => RAMDIN1(83), IN3 => 
                           RAM_12_83_port, IN4 => n5456, Q => n514);
   U511 : AO22X1 port map( IN1 => n5480, IN2 => RAMDIN1(84), IN3 => 
                           RAM_12_84_port, IN4 => n5456, Q => n515);
   U512 : AO22X1 port map( IN1 => n5480, IN2 => RAMDIN1(85), IN3 => 
                           RAM_12_85_port, IN4 => n5456, Q => n516);
   U513 : AO22X1 port map( IN1 => n5480, IN2 => RAMDIN1(86), IN3 => 
                           RAM_12_86_port, IN4 => n5456, Q => n517);
   U514 : AO22X1 port map( IN1 => n5480, IN2 => RAMDIN1(87), IN3 => 
                           RAM_12_87_port, IN4 => n5456, Q => n518);
   U515 : AO22X1 port map( IN1 => RAMDIN1(88), IN2 => n5480, IN3 => 
                           RAM_12_88_port, IN4 => n5456, Q => n519);
   U516 : AO22X1 port map( IN1 => n5481, IN2 => RAMDIN1(89), IN3 => 
                           RAM_12_89_port, IN4 => n5456, Q => n520);
   U517 : AO22X1 port map( IN1 => n5481, IN2 => RAMDIN1(90), IN3 => 
                           RAM_12_90_port, IN4 => n5456, Q => n521);
   U518 : AO22X1 port map( IN1 => n5481, IN2 => RAMDIN1(91), IN3 => 
                           RAM_12_91_port, IN4 => n5456, Q => n522);
   U519 : AO22X1 port map( IN1 => n5481, IN2 => RAMDIN1(92), IN3 => 
                           RAM_12_92_port, IN4 => n5455, Q => n523);
   U520 : AO22X1 port map( IN1 => n5481, IN2 => RAMDIN1(93), IN3 => 
                           RAM_12_93_port, IN4 => n5455, Q => n524);
   U521 : AO22X1 port map( IN1 => n5482, IN2 => RAMDIN1(94), IN3 => 
                           RAM_12_94_port, IN4 => n5455, Q => n525);
   U522 : AO22X1 port map( IN1 => n5482, IN2 => RAMDIN1(95), IN3 => 
                           RAM_12_95_port, IN4 => n5455, Q => n526);
   U523 : AO22X1 port map( IN1 => n5482, IN2 => RAMDIN1(96), IN3 => 
                           RAM_12_96_port, IN4 => n5455, Q => n527);
   U524 : AO22X1 port map( IN1 => n5482, IN2 => RAMDIN1(97), IN3 => 
                           RAM_12_97_port, IN4 => n5455, Q => n528);
   U525 : AO22X1 port map( IN1 => n5482, IN2 => RAMDIN1(98), IN3 => 
                           RAM_12_98_port, IN4 => n5455, Q => n529);
   U526 : AO22X1 port map( IN1 => n5483, IN2 => n2502, IN3 => RAM_12_99_port, 
                           IN4 => n5455, Q => n530);
   U527 : AO22X1 port map( IN1 => n5483, IN2 => RAMDIN1(100), IN3 => 
                           RAM_12_100_port, IN4 => n5455, Q => n531);
   U528 : AO22X1 port map( IN1 => n5483, IN2 => RAMDIN1(101), IN3 => 
                           RAM_12_101_port, IN4 => n5455, Q => n532);
   U529 : AO22X1 port map( IN1 => n5483, IN2 => RAMDIN1(102), IN3 => 
                           RAM_12_102_port, IN4 => n5455, Q => n533);
   U530 : AO22X1 port map( IN1 => n5483, IN2 => RAMDIN1(103), IN3 => 
                           RAM_12_103_port, IN4 => n5455, Q => n534);
   U531 : AO22X1 port map( IN1 => n5484, IN2 => RAMDIN1(104), IN3 => 
                           RAM_12_104_port, IN4 => n5454, Q => n535);
   U532 : AO22X1 port map( IN1 => n5484, IN2 => RAMDIN1(105), IN3 => 
                           RAM_12_105_port, IN4 => n5454, Q => n536);
   U533 : AO22X1 port map( IN1 => n5484, IN2 => RAMDIN1(106), IN3 => 
                           RAM_12_106_port, IN4 => n5454, Q => n537);
   U534 : AO22X1 port map( IN1 => n5484, IN2 => RAMDIN1(107), IN3 => 
                           RAM_12_107_port, IN4 => n5454, Q => n538);
   U535 : AO22X1 port map( IN1 => n5484, IN2 => RAMDIN1(108), IN3 => 
                           RAM_12_108_port, IN4 => n5454, Q => n539);
   U536 : AO22X1 port map( IN1 => n5485, IN2 => RAMDIN1(109), IN3 => 
                           RAM_12_109_port, IN4 => n5454, Q => n540);
   U537 : AO22X1 port map( IN1 => RAMDIN1(110), IN2 => n5485, IN3 => 
                           RAM_12_110_port, IN4 => n5454, Q => n541);
   U538 : AO22X1 port map( IN1 => n5485, IN2 => RAMDIN1(111), IN3 => 
                           RAM_12_111_port, IN4 => n5454, Q => n542);
   U539 : AO22X1 port map( IN1 => RAMDIN1(112), IN2 => n5485, IN3 => 
                           RAM_12_112_port, IN4 => n5454, Q => n543);
   U540 : AO22X1 port map( IN1 => n5485, IN2 => RAMDIN1(113), IN3 => 
                           RAM_12_113_port, IN4 => n5454, Q => n544);
   U541 : AO22X1 port map( IN1 => n5486, IN2 => RAMDIN1(114), IN3 => 
                           RAM_12_114_port, IN4 => n5454, Q => n545);
   U542 : AO22X1 port map( IN1 => n5486, IN2 => RAMDIN1(115), IN3 => 
                           RAM_12_115_port, IN4 => n5454, Q => n546);
   U543 : AO22X1 port map( IN1 => n5486, IN2 => RAMDIN1(116), IN3 => 
                           RAM_12_116_port, IN4 => n5453, Q => n547);
   U544 : AO22X1 port map( IN1 => n5486, IN2 => RAMDIN1(117), IN3 => 
                           RAM_12_117_port, IN4 => n5453, Q => n548);
   U545 : AO22X1 port map( IN1 => n5486, IN2 => RAMDIN1(118), IN3 => 
                           RAM_12_118_port, IN4 => n5453, Q => n549);
   U546 : AO22X1 port map( IN1 => n5487, IN2 => RAMDIN1(119), IN3 => 
                           RAM_12_119_port, IN4 => n5453, Q => n550);
   U547 : AO22X1 port map( IN1 => n5487, IN2 => RAMDIN1(120), IN3 => 
                           RAM_12_120_port, IN4 => n5453, Q => n551);
   U548 : AO22X1 port map( IN1 => n5487, IN2 => RAMDIN1(121), IN3 => 
                           RAM_12_121_port, IN4 => n5453, Q => n552);
   U549 : AO22X1 port map( IN1 => n5487, IN2 => RAMDIN1(122), IN3 => 
                           RAM_12_122_port, IN4 => n5453, Q => n553);
   U550 : AO22X1 port map( IN1 => n5487, IN2 => RAMDIN1(123), IN3 => 
                           RAM_12_123_port, IN4 => n5453, Q => n554);
   U551 : AO22X1 port map( IN1 => n5488, IN2 => RAMDIN1(124), IN3 => 
                           RAM_12_124_port, IN4 => n5453, Q => n555);
   U552 : AO22X1 port map( IN1 => n5488, IN2 => RAMDIN1(125), IN3 => 
                           RAM_12_125_port, IN4 => n5453, Q => n556);
   U553 : AO22X1 port map( IN1 => n5488, IN2 => RAMDIN1(126), IN3 => 
                           RAM_12_126_port, IN4 => n5453, Q => n557);
   U554 : AO22X1 port map( IN1 => RAMDIN1(127), IN2 => n5488, IN3 => 
                           RAM_12_127_port, IN4 => n5453, Q => n558);
   U555 : AO22X1 port map( IN1 => n5426, IN2 => RAMDIN1(0), IN3 => 
                           RAM_11_0_port, IN4 => n5422, Q => n559);
   U556 : AO22X1 port map( IN1 => n5425, IN2 => RAMDIN1(1), IN3 => 
                           RAM_11_1_port, IN4 => n5422, Q => n560);
   U557 : AO22X1 port map( IN1 => n5424, IN2 => RAMDIN1(2), IN3 => 
                           RAM_11_2_port, IN4 => n5422, Q => n561);
   U558 : AO22X1 port map( IN1 => n5424, IN2 => RAMDIN1(3), IN3 => 
                           RAM_11_3_port, IN4 => n5422, Q => n562);
   U559 : AO22X1 port map( IN1 => n5444, IN2 => RAMDIN1(4), IN3 => 
                           RAM_11_4_port, IN4 => n5422, Q => n563);
   U560 : AO22X1 port map( IN1 => n5446, IN2 => RAMDIN1(5), IN3 => 
                           RAM_11_5_port, IN4 => n5422, Q => n564);
   U561 : AO22X1 port map( IN1 => n5445, IN2 => RAMDIN1(6), IN3 => 
                           RAM_11_6_port, IN4 => n5422, Q => n565);
   U562 : AO22X1 port map( IN1 => n5444, IN2 => RAMDIN1(7), IN3 => 
                           RAM_11_7_port, IN4 => n5422, Q => n566);
   U563 : AO22X1 port map( IN1 => n5446, IN2 => RAMDIN1(8), IN3 => 
                           RAM_11_8_port, IN4 => n5421, Q => n567);
   U564 : AO22X1 port map( IN1 => n5446, IN2 => RAMDIN1(9), IN3 => 
                           RAM_11_9_port, IN4 => n5421, Q => n568);
   U565 : AO22X1 port map( IN1 => n5445, IN2 => RAMDIN1(10), IN3 => 
                           RAM_11_10_port, IN4 => n5421, Q => n569);
   U566 : AO22X1 port map( IN1 => n5444, IN2 => RAMDIN1(11), IN3 => 
                           RAM_11_11_port, IN4 => n5421, Q => n570);
   U567 : AO22X1 port map( IN1 => n5446, IN2 => RAMDIN1(12), IN3 => 
                           RAM_11_12_port, IN4 => n5421, Q => n571);
   U568 : AO22X1 port map( IN1 => n5445, IN2 => RAMDIN1(13), IN3 => 
                           RAM_11_13_port, IN4 => n5421, Q => n572);
   U569 : AO22X1 port map( IN1 => RAMDIN1(14), IN2 => n5425, IN3 => 
                           RAM_11_14_port, IN4 => n5421, Q => n573);
   U570 : AO22X1 port map( IN1 => n5425, IN2 => RAMDIN1(15), IN3 => 
                           RAM_11_15_port, IN4 => n5421, Q => n574);
   U571 : AO22X1 port map( IN1 => RAMDIN1(16), IN2 => n5425, IN3 => 
                           RAM_11_16_port, IN4 => n5421, Q => n575);
   U572 : AO22X1 port map( IN1 => n5425, IN2 => RAMDIN1(17), IN3 => 
                           RAM_11_17_port, IN4 => n5421, Q => n576);
   U573 : AO22X1 port map( IN1 => n5425, IN2 => RAMDIN1(18), IN3 => 
                           RAM_11_18_port, IN4 => n5421, Q => n577);
   U574 : AO22X1 port map( IN1 => n5426, IN2 => RAMDIN1(19), IN3 => 
                           RAM_11_19_port, IN4 => n5421, Q => n578);
   U575 : AO22X1 port map( IN1 => n5426, IN2 => RAMDIN1(20), IN3 => 
                           RAM_11_20_port, IN4 => n5420, Q => n579);
   U576 : AO22X1 port map( IN1 => n5426, IN2 => RAMDIN1(21), IN3 => 
                           RAM_11_21_port, IN4 => n5420, Q => n580);
   U577 : AO22X1 port map( IN1 => n5426, IN2 => n2249, IN3 => RAM_11_22_port, 
                           IN4 => n5420, Q => n581);
   U578 : AO22X1 port map( IN1 => n5426, IN2 => RAMDIN1(23), IN3 => 
                           RAM_11_23_port, IN4 => n5420, Q => n582);
   U579 : AO22X1 port map( IN1 => n5427, IN2 => n2106, IN3 => RAM_11_24_port, 
                           IN4 => n5420, Q => n583);
   U580 : AO22X1 port map( IN1 => n5427, IN2 => RAMDIN1(25), IN3 => 
                           RAM_11_25_port, IN4 => n5420, Q => n584);
   U581 : AO22X1 port map( IN1 => n5427, IN2 => RAMDIN1(26), IN3 => 
                           RAM_11_26_port, IN4 => n5420, Q => n585);
   U582 : AO22X1 port map( IN1 => n5427, IN2 => RAMDIN1(27), IN3 => 
                           RAM_11_27_port, IN4 => n5420, Q => n586);
   U583 : AO22X1 port map( IN1 => RAMDIN1(28), IN2 => n5427, IN3 => 
                           RAM_11_28_port, IN4 => n5420, Q => n587);
   U584 : AO22X1 port map( IN1 => n5428, IN2 => RAMDIN1(29), IN3 => 
                           RAM_11_29_port, IN4 => n5420, Q => n588);
   U585 : AO22X1 port map( IN1 => n5428, IN2 => RAMDIN1(30), IN3 => 
                           RAM_11_30_port, IN4 => n5420, Q => n589);
   U586 : AO22X1 port map( IN1 => n5428, IN2 => RAMDIN1(31), IN3 => 
                           RAM_11_31_port, IN4 => n5420, Q => n590);
   U587 : AO22X1 port map( IN1 => n5428, IN2 => RAMDIN1(32), IN3 => 
                           RAM_11_32_port, IN4 => n5419, Q => n591);
   U588 : AO22X1 port map( IN1 => n5428, IN2 => RAMDIN1(33), IN3 => 
                           RAM_11_33_port, IN4 => n5419, Q => n592);
   U589 : AO22X1 port map( IN1 => n5425, IN2 => RAMDIN1(34), IN3 => 
                           RAM_11_34_port, IN4 => n5419, Q => n593);
   U590 : AO22X1 port map( IN1 => n5427, IN2 => RAMDIN1(35), IN3 => 
                           RAM_11_35_port, IN4 => n5419, Q => n594);
   U591 : AO22X1 port map( IN1 => n5428, IN2 => RAMDIN1(36), IN3 => 
                           RAM_11_36_port, IN4 => n5419, Q => n595);
   U592 : AO22X1 port map( IN1 => n5427, IN2 => n2559, IN3 => RAM_11_37_port, 
                           IN4 => n5419, Q => n596);
   U593 : AO22X1 port map( IN1 => n5428, IN2 => RAMDIN1(38), IN3 => 
                           RAM_11_38_port, IN4 => n5419, Q => n597);
   U594 : AO22X1 port map( IN1 => n5429, IN2 => RAMDIN1(39), IN3 => 
                           RAM_11_39_port, IN4 => n5419, Q => n598);
   U595 : AO22X1 port map( IN1 => n5429, IN2 => RAMDIN1(40), IN3 => 
                           RAM_11_40_port, IN4 => n5419, Q => n599);
   U596 : AO22X1 port map( IN1 => n5429, IN2 => n2507, IN3 => RAM_11_41_port, 
                           IN4 => n5419, Q => n600);
   U597 : AO22X1 port map( IN1 => n5429, IN2 => RAMDIN1(42), IN3 => 
                           RAM_11_42_port, IN4 => n5419, Q => n601);
   U598 : AO22X1 port map( IN1 => n5429, IN2 => n2561, IN3 => RAM_11_43_port, 
                           IN4 => n5419, Q => n602);
   U599 : AO22X1 port map( IN1 => n5430, IN2 => RAMDIN1(44), IN3 => 
                           RAM_11_44_port, IN4 => n5418, Q => n603);
   U600 : AO22X1 port map( IN1 => n5430, IN2 => RAMDIN1(45), IN3 => 
                           RAM_11_45_port, IN4 => n5418, Q => n604);
   U601 : AO22X1 port map( IN1 => RAMDIN1(46), IN2 => n5430, IN3 => 
                           RAM_11_46_port, IN4 => n5418, Q => n605);
   U602 : AO22X1 port map( IN1 => n5430, IN2 => RAMDIN1(47), IN3 => 
                           RAM_11_47_port, IN4 => n5418, Q => n606);
   U603 : AO22X1 port map( IN1 => n5430, IN2 => n2557, IN3 => RAM_11_48_port, 
                           IN4 => n5418, Q => n607);
   U604 : AO22X1 port map( IN1 => n5431, IN2 => RAMDIN1(49), IN3 => 
                           RAM_11_49_port, IN4 => n5418, Q => n608);
   U605 : AO22X1 port map( IN1 => n5431, IN2 => RAMDIN1(50), IN3 => 
                           RAM_11_50_port, IN4 => n5418, Q => n609);
   U606 : AO22X1 port map( IN1 => n5431, IN2 => RAMDIN1(51), IN3 => 
                           RAM_11_51_port, IN4 => n5418, Q => n610);
   U607 : AO22X1 port map( IN1 => n5431, IN2 => n2, IN3 => RAM_11_52_port, IN4 
                           => n5418, Q => n611);
   U608 : AO22X1 port map( IN1 => n5431, IN2 => RAMDIN1(53), IN3 => 
                           RAM_11_53_port, IN4 => n5418, Q => n612);
   U609 : AO22X1 port map( IN1 => n5432, IN2 => RAMDIN1(54), IN3 => 
                           RAM_11_54_port, IN4 => n5418, Q => n613);
   U610 : AO22X1 port map( IN1 => n5432, IN2 => RAMDIN1(55), IN3 => 
                           RAM_11_55_port, IN4 => n5418, Q => n614);
   U611 : AO22X1 port map( IN1 => n5432, IN2 => RAMDIN1(56), IN3 => 
                           RAM_11_56_port, IN4 => n5417, Q => n615);
   U612 : AO22X1 port map( IN1 => RAMDIN1(57), IN2 => n5432, IN3 => 
                           RAM_11_57_port, IN4 => n5417, Q => n616);
   U613 : AO22X1 port map( IN1 => n5432, IN2 => RAMDIN1(58), IN3 => 
                           RAM_11_58_port, IN4 => n5417, Q => n617);
   U614 : AO22X1 port map( IN1 => n5433, IN2 => RAMDIN1(59), IN3 => 
                           RAM_11_59_port, IN4 => n5417, Q => n618);
   U615 : AO22X1 port map( IN1 => n5433, IN2 => RAMDIN1(60), IN3 => 
                           RAM_11_60_port, IN4 => n5417, Q => n619);
   U616 : AO22X1 port map( IN1 => n5433, IN2 => RAMDIN1(61), IN3 => 
                           RAM_11_61_port, IN4 => n5417, Q => n620);
   U617 : AO22X1 port map( IN1 => n5433, IN2 => RAMDIN1(62), IN3 => 
                           RAM_11_62_port, IN4 => n5417, Q => n621);
   U618 : AO22X1 port map( IN1 => n5433, IN2 => RAMDIN1(63), IN3 => 
                           RAM_11_63_port, IN4 => n5417, Q => n622);
   U619 : AO22X1 port map( IN1 => n5434, IN2 => RAMDIN1(64), IN3 => 
                           RAM_11_64_port, IN4 => n5417, Q => n623);
   U620 : AO22X1 port map( IN1 => n5434, IN2 => RAMDIN1(65), IN3 => 
                           RAM_11_65_port, IN4 => n5417, Q => n624);
   U621 : AO22X1 port map( IN1 => RAMDIN1(66), IN2 => n5434, IN3 => 
                           RAM_11_66_port, IN4 => n5417, Q => n625);
   U622 : AO22X1 port map( IN1 => n5434, IN2 => RAMDIN1(67), IN3 => 
                           RAM_11_67_port, IN4 => n5417, Q => n626);
   U623 : AO22X1 port map( IN1 => n5434, IN2 => RAMDIN1(68), IN3 => 
                           RAM_11_68_port, IN4 => n5416, Q => n627);
   U624 : AO22X1 port map( IN1 => n5435, IN2 => RAMDIN1(69), IN3 => 
                           RAM_11_69_port, IN4 => n5416, Q => n628);
   U625 : AO22X1 port map( IN1 => n5435, IN2 => RAMDIN1(70), IN3 => 
                           RAM_11_70_port, IN4 => n5416, Q => n629);
   U626 : AO22X1 port map( IN1 => n5435, IN2 => RAMDIN1(71), IN3 => 
                           RAM_11_71_port, IN4 => n5416, Q => n630);
   U627 : AO22X1 port map( IN1 => n5435, IN2 => RAMDIN1(72), IN3 => 
                           RAM_11_72_port, IN4 => n5416, Q => n631);
   U628 : AO22X1 port map( IN1 => n5435, IN2 => RAMDIN1(73), IN3 => 
                           RAM_11_73_port, IN4 => n5416, Q => n632);
   U629 : AO22X1 port map( IN1 => n5436, IN2 => RAMDIN1(74), IN3 => 
                           RAM_11_74_port, IN4 => n5416, Q => n633);
   U630 : AO22X1 port map( IN1 => n5436, IN2 => RAMDIN1(75), IN3 => 
                           RAM_11_75_port, IN4 => n5416, Q => n634);
   U631 : AO22X1 port map( IN1 => n5436, IN2 => RAMDIN1(76), IN3 => 
                           RAM_11_76_port, IN4 => n5416, Q => n635);
   U632 : AO22X1 port map( IN1 => n5436, IN2 => RAMDIN1(77), IN3 => 
                           RAM_11_77_port, IN4 => n5416, Q => n636);
   U633 : AO22X1 port map( IN1 => n5436, IN2 => RAMDIN1(78), IN3 => 
                           RAM_11_78_port, IN4 => n5416, Q => n637);
   U634 : AO22X1 port map( IN1 => n5437, IN2 => RAMDIN1(79), IN3 => 
                           RAM_11_79_port, IN4 => n5416, Q => n638);
   U635 : AO22X1 port map( IN1 => RAMDIN1(80), IN2 => n5437, IN3 => 
                           RAM_11_80_port, IN4 => n5415, Q => n639);
   U636 : AO22X1 port map( IN1 => n5437, IN2 => RAMDIN1(81), IN3 => 
                           RAM_11_81_port, IN4 => n5415, Q => n640);
   U637 : AO22X1 port map( IN1 => n5437, IN2 => RAMDIN1(82), IN3 => 
                           RAM_11_82_port, IN4 => n5415, Q => n641);
   U638 : AO22X1 port map( IN1 => RAMDIN1(83), IN2 => n5437, IN3 => 
                           RAM_11_83_port, IN4 => n5415, Q => n642);
   U639 : AO22X1 port map( IN1 => n5438, IN2 => RAMDIN1(84), IN3 => 
                           RAM_11_84_port, IN4 => n5415, Q => n643);
   U640 : AO22X1 port map( IN1 => n5438, IN2 => RAMDIN1(85), IN3 => 
                           RAM_11_85_port, IN4 => n5415, Q => n644);
   U641 : AO22X1 port map( IN1 => n5438, IN2 => RAMDIN1(86), IN3 => 
                           RAM_11_86_port, IN4 => n5415, Q => n645);
   U642 : AO22X1 port map( IN1 => n5438, IN2 => RAMDIN1(87), IN3 => 
                           RAM_11_87_port, IN4 => n5415, Q => n646);
   U643 : AO22X1 port map( IN1 => RAMDIN1(88), IN2 => n5438, IN3 => 
                           RAM_11_88_port, IN4 => n5415, Q => n647);
   U644 : AO22X1 port map( IN1 => n5439, IN2 => RAMDIN1(89), IN3 => 
                           RAM_11_89_port, IN4 => n5415, Q => n648);
   U645 : AO22X1 port map( IN1 => n5439, IN2 => RAMDIN1(90), IN3 => 
                           RAM_11_90_port, IN4 => n5415, Q => n649);
   U646 : AO22X1 port map( IN1 => RAMDIN1(91), IN2 => n5439, IN3 => 
                           RAM_11_91_port, IN4 => n5415, Q => n650);
   U647 : AO22X1 port map( IN1 => n5439, IN2 => RAMDIN1(92), IN3 => 
                           RAM_11_92_port, IN4 => n5414, Q => n651);
   U648 : AO22X1 port map( IN1 => n5439, IN2 => RAMDIN1(93), IN3 => 
                           RAM_11_93_port, IN4 => n5414, Q => n652);
   U649 : AO22X1 port map( IN1 => n5440, IN2 => RAMDIN1(94), IN3 => 
                           RAM_11_94_port, IN4 => n5414, Q => n653);
   U650 : AO22X1 port map( IN1 => n5440, IN2 => RAMDIN1(95), IN3 => 
                           RAM_11_95_port, IN4 => n5414, Q => n654);
   U651 : AO22X1 port map( IN1 => n5440, IN2 => RAMDIN1(96), IN3 => 
                           RAM_11_96_port, IN4 => n5414, Q => n655);
   U652 : AO22X1 port map( IN1 => n5440, IN2 => RAMDIN1(97), IN3 => 
                           RAM_11_97_port, IN4 => n5414, Q => n656);
   U653 : AO22X1 port map( IN1 => n5440, IN2 => RAMDIN1(98), IN3 => 
                           RAM_11_98_port, IN4 => n5414, Q => n657);
   U654 : AO22X1 port map( IN1 => n5441, IN2 => n2102, IN3 => RAM_11_99_port, 
                           IN4 => n5414, Q => n658);
   U655 : AO22X1 port map( IN1 => n5441, IN2 => RAMDIN1(100), IN3 => 
                           RAM_11_100_port, IN4 => n5414, Q => n659);
   U656 : AO22X1 port map( IN1 => n5441, IN2 => RAMDIN1(101), IN3 => 
                           RAM_11_101_port, IN4 => n5414, Q => n660);
   U657 : AO22X1 port map( IN1 => n5441, IN2 => RAMDIN1(102), IN3 => 
                           RAM_11_102_port, IN4 => n5414, Q => n661);
   U658 : AO22X1 port map( IN1 => n5441, IN2 => RAMDIN1(103), IN3 => 
                           RAM_11_103_port, IN4 => n5414, Q => n662);
   U659 : AO22X1 port map( IN1 => n5442, IN2 => RAMDIN1(104), IN3 => 
                           RAM_11_104_port, IN4 => n5413, Q => n663);
   U660 : AO22X1 port map( IN1 => n5442, IN2 => RAMDIN1(105), IN3 => 
                           RAM_11_105_port, IN4 => n5413, Q => n664);
   U661 : AO22X1 port map( IN1 => n5442, IN2 => RAMDIN1(106), IN3 => 
                           RAM_11_106_port, IN4 => n5413, Q => n665);
   U662 : AO22X1 port map( IN1 => n5442, IN2 => RAMDIN1(107), IN3 => 
                           RAM_11_107_port, IN4 => n5413, Q => n666);
   U663 : AO22X1 port map( IN1 => n5442, IN2 => RAMDIN1(108), IN3 => 
                           RAM_11_108_port, IN4 => n5413, Q => n667);
   U664 : AO22X1 port map( IN1 => n5443, IN2 => RAMDIN1(109), IN3 => 
                           RAM_11_109_port, IN4 => n5413, Q => n668);
   U665 : AO22X1 port map( IN1 => RAMDIN1(110), IN2 => n5443, IN3 => 
                           RAM_11_110_port, IN4 => n5413, Q => n669);
   U666 : AO22X1 port map( IN1 => n5443, IN2 => RAMDIN1(111), IN3 => 
                           RAM_11_111_port, IN4 => n5413, Q => n670);
   U667 : AO22X1 port map( IN1 => RAMDIN1(112), IN2 => n5443, IN3 => 
                           RAM_11_112_port, IN4 => n5413, Q => n671);
   U668 : AO22X1 port map( IN1 => n5443, IN2 => RAMDIN1(113), IN3 => 
                           RAM_11_113_port, IN4 => n5413, Q => n672);
   U669 : AO22X1 port map( IN1 => n5444, IN2 => RAMDIN1(114), IN3 => 
                           RAM_11_114_port, IN4 => n5413, Q => n673);
   U670 : AO22X1 port map( IN1 => n5444, IN2 => RAMDIN1(115), IN3 => 
                           RAM_11_115_port, IN4 => n5413, Q => n674);
   U671 : AO22X1 port map( IN1 => n5444, IN2 => RAMDIN1(116), IN3 => 
                           RAM_11_116_port, IN4 => n5412, Q => n675);
   U672 : AO22X1 port map( IN1 => n5444, IN2 => RAMDIN1(117), IN3 => 
                           RAM_11_117_port, IN4 => n5412, Q => n676);
   U673 : AO22X1 port map( IN1 => n5444, IN2 => RAMDIN1(118), IN3 => 
                           RAM_11_118_port, IN4 => n5412, Q => n677);
   U674 : AO22X1 port map( IN1 => n5445, IN2 => RAMDIN1(119), IN3 => 
                           RAM_11_119_port, IN4 => n5412, Q => n678);
   U675 : AO22X1 port map( IN1 => n5445, IN2 => RAMDIN1(120), IN3 => 
                           RAM_11_120_port, IN4 => n5412, Q => n679);
   U676 : AO22X1 port map( IN1 => n5445, IN2 => RAMDIN1(121), IN3 => 
                           RAM_11_121_port, IN4 => n5412, Q => n680);
   U677 : AO22X1 port map( IN1 => RAMDIN1(122), IN2 => n5445, IN3 => 
                           RAM_11_122_port, IN4 => n5412, Q => n681);
   U678 : AO22X1 port map( IN1 => n5445, IN2 => RAMDIN1(123), IN3 => 
                           RAM_11_123_port, IN4 => n5412, Q => n682);
   U679 : AO22X1 port map( IN1 => n5446, IN2 => RAMDIN1(124), IN3 => 
                           RAM_11_124_port, IN4 => n5412, Q => n683);
   U680 : AO22X1 port map( IN1 => n5446, IN2 => RAMDIN1(125), IN3 => 
                           RAM_11_125_port, IN4 => n5412, Q => n684);
   U681 : AO22X1 port map( IN1 => n5446, IN2 => RAMDIN1(126), IN3 => 
                           RAM_11_126_port, IN4 => n5412, Q => n685);
   U682 : AO22X1 port map( IN1 => RAMDIN1(127), IN2 => n5446, IN3 => 
                           RAM_11_127_port, IN4 => n5412, Q => n686);
   U683 : AO22X1 port map( IN1 => n5386, IN2 => RAMDIN1(0), IN3 => 
                           RAM_10_0_port, IN4 => n5381, Q => n687);
   U684 : AO22X1 port map( IN1 => n5384, IN2 => RAMDIN1(1), IN3 => 
                           RAM_10_1_port, IN4 => n5381, Q => n688);
   U685 : AO22X1 port map( IN1 => n5382, IN2 => RAMDIN1(2), IN3 => 
                           RAM_10_2_port, IN4 => n5381, Q => n689);
   U686 : AO22X1 port map( IN1 => n5382, IN2 => RAMDIN1(3), IN3 => 
                           RAM_10_3_port, IN4 => n5381, Q => n690);
   U687 : AO22X1 port map( IN1 => n5403, IN2 => RAMDIN1(4), IN3 => 
                           RAM_10_4_port, IN4 => n5381, Q => n691);
   U688 : AO22X1 port map( IN1 => n5405, IN2 => RAMDIN1(5), IN3 => 
                           RAM_10_5_port, IN4 => n5381, Q => n692);
   U689 : AO22X1 port map( IN1 => n5404, IN2 => RAMDIN1(6), IN3 => 
                           RAM_10_6_port, IN4 => n5381, Q => n693);
   U690 : AO22X1 port map( IN1 => n5403, IN2 => RAMDIN1(7), IN3 => 
                           RAM_10_7_port, IN4 => n5381, Q => n694);
   U691 : AO22X1 port map( IN1 => n5405, IN2 => RAMDIN1(8), IN3 => 
                           RAM_10_8_port, IN4 => n5380, Q => n695);
   U692 : AO22X1 port map( IN1 => n5405, IN2 => RAMDIN1(9), IN3 => 
                           RAM_10_9_port, IN4 => n5380, Q => n696);
   U693 : AO22X1 port map( IN1 => n5404, IN2 => RAMDIN1(10), IN3 => 
                           RAM_10_10_port, IN4 => n5380, Q => n697);
   U694 : AO22X1 port map( IN1 => n5403, IN2 => RAMDIN1(11), IN3 => 
                           RAM_10_11_port, IN4 => n5380, Q => n698);
   U695 : AO22X1 port map( IN1 => n5405, IN2 => RAMDIN1(12), IN3 => 
                           RAM_10_12_port, IN4 => n5380, Q => n699);
   U696 : AO22X1 port map( IN1 => n5404, IN2 => RAMDIN1(13), IN3 => 
                           RAM_10_13_port, IN4 => n5380, Q => n700);
   U697 : AO22X1 port map( IN1 => RAMDIN1(14), IN2 => n5384, IN3 => 
                           RAM_10_14_port, IN4 => n5380, Q => n701);
   U698 : AO22X1 port map( IN1 => n5384, IN2 => RAMDIN1(15), IN3 => 
                           RAM_10_15_port, IN4 => n5380, Q => n702);
   U699 : AO22X1 port map( IN1 => RAMDIN1(16), IN2 => n5384, IN3 => 
                           RAM_10_16_port, IN4 => n5380, Q => n703);
   U700 : AO22X1 port map( IN1 => n5384, IN2 => RAMDIN1(17), IN3 => 
                           RAM_10_17_port, IN4 => n5380, Q => n704);
   U701 : AO22X1 port map( IN1 => n5384, IN2 => RAMDIN1(18), IN3 => 
                           RAM_10_18_port, IN4 => n5380, Q => n705);
   U702 : AO22X1 port map( IN1 => n5386, IN2 => RAMDIN1(19), IN3 => 
                           RAM_10_19_port, IN4 => n5380, Q => n706);
   U703 : AO22X1 port map( IN1 => n5385, IN2 => RAMDIN1(20), IN3 => 
                           RAM_10_20_port, IN4 => n5379, Q => n707);
   U704 : AO22X1 port map( IN1 => n5385, IN2 => RAMDIN1(21), IN3 => 
                           RAM_10_21_port, IN4 => n5379, Q => n708);
   U705 : AO22X1 port map( IN1 => n5384, IN2 => n2249, IN3 => RAM_10_22_port, 
                           IN4 => n5379, Q => n709);
   U706 : AO22X1 port map( IN1 => n5387, IN2 => RAMDIN1(23), IN3 => 
                           RAM_10_23_port, IN4 => n5379, Q => n710);
   U707 : AO22X1 port map( IN1 => n5385, IN2 => n2106, IN3 => RAM_10_24_port, 
                           IN4 => n5379, Q => n711);
   U708 : AO22X1 port map( IN1 => n5385, IN2 => RAMDIN1(25), IN3 => 
                           RAM_10_25_port, IN4 => n5379, Q => n712);
   U709 : AO22X1 port map( IN1 => n5385, IN2 => RAMDIN1(26), IN3 => 
                           RAM_10_26_port, IN4 => n5379, Q => n713);
   U710 : AO22X1 port map( IN1 => n5385, IN2 => RAMDIN1(27), IN3 => 
                           RAM_10_27_port, IN4 => n5379, Q => n714);
   U711 : AO22X1 port map( IN1 => RAMDIN1(28), IN2 => n5385, IN3 => 
                           RAM_10_28_port, IN4 => n5379, Q => n715);
   U712 : AO22X1 port map( IN1 => n5386, IN2 => RAMDIN1(29), IN3 => 
                           RAM_10_29_port, IN4 => n5379, Q => n716);
   U713 : AO22X1 port map( IN1 => RAMDIN1(30), IN2 => n5386, IN3 => 
                           RAM_10_30_port, IN4 => n5379, Q => n717);
   U714 : AO22X1 port map( IN1 => n5386, IN2 => RAMDIN1(31), IN3 => 
                           RAM_10_31_port, IN4 => n5379, Q => n718);
   U715 : AO22X1 port map( IN1 => n5386, IN2 => RAMDIN1(32), IN3 => 
                           RAM_10_32_port, IN4 => n5378, Q => n719);
   U716 : AO22X1 port map( IN1 => n5386, IN2 => RAMDIN1(33), IN3 => 
                           RAM_10_33_port, IN4 => n5378, Q => n720);
   U717 : AO22X1 port map( IN1 => n5387, IN2 => RAMDIN1(34), IN3 => 
                           RAM_10_34_port, IN4 => n5378, Q => n721);
   U718 : AO22X1 port map( IN1 => n5387, IN2 => RAMDIN1(35), IN3 => 
                           RAM_10_35_port, IN4 => n5378, Q => n722);
   U719 : AO22X1 port map( IN1 => n5387, IN2 => RAMDIN1(36), IN3 => 
                           RAM_10_36_port, IN4 => n5378, Q => n723);
   U720 : AO22X1 port map( IN1 => n5387, IN2 => n2558, IN3 => RAM_10_37_port, 
                           IN4 => n5378, Q => n724);
   U721 : AO22X1 port map( IN1 => n5387, IN2 => RAMDIN1(38), IN3 => 
                           RAM_10_38_port, IN4 => n5378, Q => n725);
   U722 : AO22X1 port map( IN1 => n5388, IN2 => RAMDIN1(39), IN3 => 
                           RAM_10_39_port, IN4 => n5378, Q => n726);
   U723 : AO22X1 port map( IN1 => n5388, IN2 => RAMDIN1(40), IN3 => 
                           RAM_10_40_port, IN4 => n5378, Q => n727);
   U724 : AO22X1 port map( IN1 => n5388, IN2 => n2104, IN3 => RAM_10_41_port, 
                           IN4 => n5378, Q => n728);
   U725 : AO22X1 port map( IN1 => n5388, IN2 => RAMDIN1(42), IN3 => 
                           RAM_10_42_port, IN4 => n5378, Q => n729);
   U726 : AO22X1 port map( IN1 => n5388, IN2 => n2101, IN3 => RAM_10_43_port, 
                           IN4 => n5378, Q => n730);
   U727 : AO22X1 port map( IN1 => RAMDIN1(44), IN2 => n5389, IN3 => 
                           RAM_10_44_port, IN4 => n5377, Q => n731);
   U728 : AO22X1 port map( IN1 => RAMDIN1(45), IN2 => n5389, IN3 => 
                           RAM_10_45_port, IN4 => n5377, Q => n732);
   U729 : AO22X1 port map( IN1 => RAMDIN1(46), IN2 => n5389, IN3 => 
                           RAM_10_46_port, IN4 => n5377, Q => n733);
   U730 : AO22X1 port map( IN1 => n5389, IN2 => RAMDIN1(47), IN3 => 
                           RAM_10_47_port, IN4 => n5377, Q => n734);
   U731 : AO22X1 port map( IN1 => n5389, IN2 => n2126, IN3 => RAM_10_48_port, 
                           IN4 => n5377, Q => n735);
   U732 : AO22X1 port map( IN1 => n5390, IN2 => RAMDIN1(49), IN3 => 
                           RAM_10_49_port, IN4 => n5377, Q => n736);
   U733 : AO22X1 port map( IN1 => n5390, IN2 => RAMDIN1(50), IN3 => 
                           RAM_10_50_port, IN4 => n5377, Q => n737);
   U734 : AO22X1 port map( IN1 => n5390, IN2 => RAMDIN1(51), IN3 => 
                           RAM_10_51_port, IN4 => n5377, Q => n738);
   U735 : AO22X1 port map( IN1 => n5390, IN2 => n2556, IN3 => RAM_10_52_port, 
                           IN4 => n5377, Q => n739);
   U736 : AO22X1 port map( IN1 => n5390, IN2 => RAMDIN1(53), IN3 => 
                           RAM_10_53_port, IN4 => n5377, Q => n740);
   U737 : AO22X1 port map( IN1 => n5391, IN2 => RAMDIN1(54), IN3 => 
                           RAM_10_54_port, IN4 => n5377, Q => n741);
   U738 : AO22X1 port map( IN1 => n5391, IN2 => RAMDIN1(55), IN3 => 
                           RAM_10_55_port, IN4 => n5377, Q => n742);
   U739 : AO22X1 port map( IN1 => n5391, IN2 => RAMDIN1(56), IN3 => 
                           RAM_10_56_port, IN4 => n5376, Q => n743);
   U740 : AO22X1 port map( IN1 => n5391, IN2 => RAMDIN1(57), IN3 => 
                           RAM_10_57_port, IN4 => n5376, Q => n744);
   U741 : AO22X1 port map( IN1 => n5391, IN2 => RAMDIN1(58), IN3 => 
                           RAM_10_58_port, IN4 => n5376, Q => n745);
   U742 : AO22X1 port map( IN1 => n5392, IN2 => RAMDIN1(59), IN3 => 
                           RAM_10_59_port, IN4 => n5376, Q => n746);
   U743 : AO22X1 port map( IN1 => n5392, IN2 => RAMDIN1(60), IN3 => 
                           RAM_10_60_port, IN4 => n5376, Q => n747);
   U744 : AO22X1 port map( IN1 => n5392, IN2 => RAMDIN1(61), IN3 => 
                           RAM_10_61_port, IN4 => n5376, Q => n748);
   U745 : AO22X1 port map( IN1 => n5392, IN2 => RAMDIN1(62), IN3 => 
                           RAM_10_62_port, IN4 => n5376, Q => n749);
   U746 : AO22X1 port map( IN1 => n5392, IN2 => RAMDIN1(63), IN3 => 
                           RAM_10_63_port, IN4 => n5376, Q => n750);
   U747 : AO22X1 port map( IN1 => n5393, IN2 => RAMDIN1(64), IN3 => 
                           RAM_10_64_port, IN4 => n5376, Q => n751);
   U748 : AO22X1 port map( IN1 => n5393, IN2 => RAMDIN1(65), IN3 => 
                           RAM_10_65_port, IN4 => n5376, Q => n752);
   U749 : AO22X1 port map( IN1 => n5393, IN2 => RAMDIN1(66), IN3 => 
                           RAM_10_66_port, IN4 => n5376, Q => n753);
   U750 : AO22X1 port map( IN1 => n5393, IN2 => RAMDIN1(67), IN3 => 
                           RAM_10_67_port, IN4 => n5376, Q => n754);
   U751 : AO22X1 port map( IN1 => n5393, IN2 => RAMDIN1(68), IN3 => 
                           RAM_10_68_port, IN4 => n5375, Q => n755);
   U752 : AO22X1 port map( IN1 => n5394, IN2 => RAMDIN1(69), IN3 => 
                           RAM_10_69_port, IN4 => n5375, Q => n756);
   U753 : AO22X1 port map( IN1 => n5394, IN2 => RAMDIN1(70), IN3 => 
                           RAM_10_70_port, IN4 => n5375, Q => n757);
   U754 : AO22X1 port map( IN1 => n5394, IN2 => RAMDIN1(71), IN3 => 
                           RAM_10_71_port, IN4 => n5375, Q => n758);
   U755 : AO22X1 port map( IN1 => n5394, IN2 => RAMDIN1(72), IN3 => 
                           RAM_10_72_port, IN4 => n5375, Q => n759);
   U756 : AO22X1 port map( IN1 => n5394, IN2 => RAMDIN1(73), IN3 => 
                           RAM_10_73_port, IN4 => n5375, Q => n760);
   U757 : AO22X1 port map( IN1 => n5395, IN2 => RAMDIN1(74), IN3 => 
                           RAM_10_74_port, IN4 => n5375, Q => n761);
   U758 : AO22X1 port map( IN1 => n5395, IN2 => RAMDIN1(75), IN3 => 
                           RAM_10_75_port, IN4 => n5375, Q => n762);
   U759 : AO22X1 port map( IN1 => n5395, IN2 => RAMDIN1(76), IN3 => 
                           RAM_10_76_port, IN4 => n5375, Q => n763);
   U760 : AO22X1 port map( IN1 => n5395, IN2 => RAMDIN1(77), IN3 => 
                           RAM_10_77_port, IN4 => n5375, Q => n764);
   U761 : AO22X1 port map( IN1 => n5395, IN2 => RAMDIN1(78), IN3 => 
                           RAM_10_78_port, IN4 => n5375, Q => n765);
   U762 : AO22X1 port map( IN1 => n5396, IN2 => RAMDIN1(79), IN3 => 
                           RAM_10_79_port, IN4 => n5375, Q => n766);
   U763 : AO22X1 port map( IN1 => RAMDIN1(80), IN2 => n5396, IN3 => 
                           RAM_10_80_port, IN4 => n5374, Q => n767);
   U764 : AO22X1 port map( IN1 => n5396, IN2 => RAMDIN1(81), IN3 => 
                           RAM_10_81_port, IN4 => n5374, Q => n768);
   U765 : AO22X1 port map( IN1 => n5396, IN2 => RAMDIN1(82), IN3 => 
                           RAM_10_82_port, IN4 => n5374, Q => n769);
   U766 : AO22X1 port map( IN1 => n5396, IN2 => RAMDIN1(83), IN3 => 
                           RAM_10_83_port, IN4 => n5374, Q => n770);
   U767 : AO22X1 port map( IN1 => n5397, IN2 => RAMDIN1(84), IN3 => 
                           RAM_10_84_port, IN4 => n5374, Q => n771);
   U768 : AO22X1 port map( IN1 => n5397, IN2 => RAMDIN1(85), IN3 => 
                           RAM_10_85_port, IN4 => n5374, Q => n772);
   U769 : AO22X1 port map( IN1 => n5397, IN2 => RAMDIN1(86), IN3 => 
                           RAM_10_86_port, IN4 => n5374, Q => n773);
   U770 : AO22X1 port map( IN1 => n5397, IN2 => RAMDIN1(87), IN3 => 
                           RAM_10_87_port, IN4 => n5374, Q => n774);
   U771 : AO22X1 port map( IN1 => RAMDIN1(88), IN2 => n5397, IN3 => 
                           RAM_10_88_port, IN4 => n5374, Q => n775);
   U772 : AO22X1 port map( IN1 => n5398, IN2 => RAMDIN1(89), IN3 => 
                           RAM_10_89_port, IN4 => n5374, Q => n776);
   U773 : AO22X1 port map( IN1 => n5398, IN2 => RAMDIN1(90), IN3 => 
                           RAM_10_90_port, IN4 => n5374, Q => n777);
   U774 : AO22X1 port map( IN1 => n5398, IN2 => RAMDIN1(91), IN3 => 
                           RAM_10_91_port, IN4 => n5374, Q => n778);
   U775 : AO22X1 port map( IN1 => n5398, IN2 => RAMDIN1(92), IN3 => 
                           RAM_10_92_port, IN4 => n5373, Q => n779);
   U776 : AO22X1 port map( IN1 => n5398, IN2 => RAMDIN1(93), IN3 => 
                           RAM_10_93_port, IN4 => n5373, Q => n780);
   U777 : AO22X1 port map( IN1 => n5399, IN2 => RAMDIN1(94), IN3 => 
                           RAM_10_94_port, IN4 => n5373, Q => n781);
   U778 : AO22X1 port map( IN1 => n5399, IN2 => RAMDIN1(95), IN3 => 
                           RAM_10_95_port, IN4 => n5373, Q => n782);
   U779 : AO22X1 port map( IN1 => n5399, IN2 => RAMDIN1(96), IN3 => 
                           RAM_10_96_port, IN4 => n5373, Q => n783);
   U780 : AO22X1 port map( IN1 => n5399, IN2 => RAMDIN1(97), IN3 => 
                           RAM_10_97_port, IN4 => n5373, Q => n784);
   U781 : AO22X1 port map( IN1 => n5399, IN2 => RAMDIN1(98), IN3 => 
                           RAM_10_98_port, IN4 => n5373, Q => n785);
   U782 : AO22X1 port map( IN1 => n5400, IN2 => n2503, IN3 => RAM_10_99_port, 
                           IN4 => n5373, Q => n786);
   U783 : AO22X1 port map( IN1 => n5400, IN2 => RAMDIN1(100), IN3 => 
                           RAM_10_100_port, IN4 => n5373, Q => n787);
   U784 : AO22X1 port map( IN1 => n5400, IN2 => RAMDIN1(101), IN3 => 
                           RAM_10_101_port, IN4 => n5373, Q => n788);
   U785 : AO22X1 port map( IN1 => n5400, IN2 => RAMDIN1(102), IN3 => 
                           RAM_10_102_port, IN4 => n5373, Q => n789);
   U786 : AO22X1 port map( IN1 => n5400, IN2 => RAMDIN1(103), IN3 => 
                           RAM_10_103_port, IN4 => n5373, Q => n790);
   U787 : AO22X1 port map( IN1 => n5401, IN2 => RAMDIN1(104), IN3 => 
                           RAM_10_104_port, IN4 => n5372, Q => n791);
   U788 : AO22X1 port map( IN1 => n5401, IN2 => RAMDIN1(105), IN3 => 
                           RAM_10_105_port, IN4 => n5372, Q => n792);
   U789 : AO22X1 port map( IN1 => n5401, IN2 => RAMDIN1(106), IN3 => 
                           RAM_10_106_port, IN4 => n5372, Q => n793);
   U790 : AO22X1 port map( IN1 => n5401, IN2 => RAMDIN1(107), IN3 => 
                           RAM_10_107_port, IN4 => n5372, Q => n794);
   U791 : AO22X1 port map( IN1 => n5401, IN2 => RAMDIN1(108), IN3 => 
                           RAM_10_108_port, IN4 => n5372, Q => n795);
   U792 : AO22X1 port map( IN1 => n5402, IN2 => RAMDIN1(109), IN3 => 
                           RAM_10_109_port, IN4 => n5372, Q => n796);
   U793 : AO22X1 port map( IN1 => RAMDIN1(110), IN2 => n5402, IN3 => 
                           RAM_10_110_port, IN4 => n5372, Q => n797);
   U794 : AO22X1 port map( IN1 => n5402, IN2 => RAMDIN1(111), IN3 => 
                           RAM_10_111_port, IN4 => n5372, Q => n798);
   U795 : AO22X1 port map( IN1 => RAMDIN1(112), IN2 => n5402, IN3 => 
                           RAM_10_112_port, IN4 => n5372, Q => n799);
   U796 : AO22X1 port map( IN1 => n5402, IN2 => RAMDIN1(113), IN3 => 
                           RAM_10_113_port, IN4 => n5372, Q => n800);
   U797 : AO22X1 port map( IN1 => n5403, IN2 => RAMDIN1(114), IN3 => 
                           RAM_10_114_port, IN4 => n5372, Q => n801);
   U798 : AO22X1 port map( IN1 => n5403, IN2 => RAMDIN1(115), IN3 => 
                           RAM_10_115_port, IN4 => n5372, Q => n802);
   U799 : AO22X1 port map( IN1 => n5403, IN2 => RAMDIN1(116), IN3 => 
                           RAM_10_116_port, IN4 => n5371, Q => n803);
   U800 : AO22X1 port map( IN1 => n5403, IN2 => RAMDIN1(117), IN3 => 
                           RAM_10_117_port, IN4 => n5371, Q => n804);
   U801 : AO22X1 port map( IN1 => n5403, IN2 => RAMDIN1(118), IN3 => 
                           RAM_10_118_port, IN4 => n5371, Q => n805);
   U802 : AO22X1 port map( IN1 => n5404, IN2 => RAMDIN1(119), IN3 => 
                           RAM_10_119_port, IN4 => n5371, Q => n806);
   U803 : AO22X1 port map( IN1 => n5404, IN2 => RAMDIN1(120), IN3 => 
                           RAM_10_120_port, IN4 => n5371, Q => n807);
   U804 : AO22X1 port map( IN1 => n5404, IN2 => RAMDIN1(121), IN3 => 
                           RAM_10_121_port, IN4 => n5371, Q => n808);
   U805 : AO22X1 port map( IN1 => n5404, IN2 => RAMDIN1(122), IN3 => 
                           RAM_10_122_port, IN4 => n5371, Q => n809);
   U806 : AO22X1 port map( IN1 => n5404, IN2 => RAMDIN1(123), IN3 => 
                           RAM_10_123_port, IN4 => n5371, Q => n810);
   U807 : AO22X1 port map( IN1 => n5405, IN2 => RAMDIN1(124), IN3 => 
                           RAM_10_124_port, IN4 => n5371, Q => n811);
   U808 : AO22X1 port map( IN1 => n5405, IN2 => RAMDIN1(125), IN3 => 
                           RAM_10_125_port, IN4 => n5371, Q => n812);
   U809 : AO22X1 port map( IN1 => n5405, IN2 => RAMDIN1(126), IN3 => 
                           RAM_10_126_port, IN4 => n5371, Q => n813);
   U810 : AO22X1 port map( IN1 => RAMDIN1(127), IN2 => n5405, IN3 => 
                           RAM_10_127_port, IN4 => n5371, Q => n814);
   U811 : AO22X1 port map( IN1 => n5343, IN2 => RAMDIN1(0), IN3 => RAM_9_0_port
                           , IN4 => n5339, Q => n815);
   U812 : AO22X1 port map( IN1 => n5342, IN2 => RAMDIN1(1), IN3 => RAM_9_1_port
                           , IN4 => n5339, Q => n816);
   U813 : AO22X1 port map( IN1 => n5341, IN2 => RAMDIN1(2), IN3 => RAM_9_2_port
                           , IN4 => n5339, Q => n817);
   U814 : AO22X1 port map( IN1 => n5341, IN2 => RAMDIN1(3), IN3 => RAM_9_3_port
                           , IN4 => n5339, Q => n818);
   U815 : AO22X1 port map( IN1 => n5362, IN2 => RAMDIN1(4), IN3 => RAM_9_4_port
                           , IN4 => n5339, Q => n819);
   U816 : AO22X1 port map( IN1 => n5364, IN2 => RAMDIN1(5), IN3 => RAM_9_5_port
                           , IN4 => n5339, Q => n820);
   U817 : AO22X1 port map( IN1 => n5363, IN2 => RAMDIN1(6), IN3 => RAM_9_6_port
                           , IN4 => n5339, Q => n821);
   U818 : AO22X1 port map( IN1 => n5362, IN2 => RAMDIN1(7), IN3 => RAM_9_7_port
                           , IN4 => n5339, Q => n822);
   U819 : AO22X1 port map( IN1 => n5364, IN2 => RAMDIN1(8), IN3 => RAM_9_8_port
                           , IN4 => n5338, Q => n823);
   U820 : AO22X1 port map( IN1 => n5364, IN2 => RAMDIN1(9), IN3 => RAM_9_9_port
                           , IN4 => n5338, Q => n824);
   U821 : AO22X1 port map( IN1 => n5363, IN2 => RAMDIN1(10), IN3 => 
                           RAM_9_10_port, IN4 => n5338, Q => n825);
   U822 : AO22X1 port map( IN1 => n5362, IN2 => RAMDIN1(11), IN3 => 
                           RAM_9_11_port, IN4 => n5338, Q => n826);
   U823 : AO22X1 port map( IN1 => n5364, IN2 => RAMDIN1(12), IN3 => 
                           RAM_9_12_port, IN4 => n5338, Q => n827);
   U824 : AO22X1 port map( IN1 => n5363, IN2 => RAMDIN1(13), IN3 => 
                           RAM_9_13_port, IN4 => n5338, Q => n828);
   U825 : AO22X1 port map( IN1 => RAMDIN1(14), IN2 => n5342, IN3 => 
                           RAM_9_14_port, IN4 => n5338, Q => n829);
   U826 : AO22X1 port map( IN1 => n5342, IN2 => RAMDIN1(15), IN3 => 
                           RAM_9_15_port, IN4 => n5338, Q => n830);
   U827 : AO22X1 port map( IN1 => RAMDIN1(16), IN2 => n5342, IN3 => 
                           RAM_9_16_port, IN4 => n5338, Q => n831);
   U828 : AO22X1 port map( IN1 => n5342, IN2 => RAMDIN1(17), IN3 => 
                           RAM_9_17_port, IN4 => n5338, Q => n832);
   U829 : AO22X1 port map( IN1 => n5342, IN2 => RAMDIN1(18), IN3 => 
                           RAM_9_18_port, IN4 => n5338, Q => n833);
   U830 : AO22X1 port map( IN1 => n5343, IN2 => RAMDIN1(19), IN3 => 
                           RAM_9_19_port, IN4 => n5338, Q => n834);
   U831 : AO22X1 port map( IN1 => n5343, IN2 => RAMDIN1(20), IN3 => 
                           RAM_9_20_port, IN4 => n5337, Q => n835);
   U832 : AO22X1 port map( IN1 => n5343, IN2 => RAMDIN1(21), IN3 => 
                           RAM_9_21_port, IN4 => n5337, Q => n836);
   U833 : AO22X1 port map( IN1 => n5343, IN2 => n2103, IN3 => RAM_9_22_port, 
                           IN4 => n5337, Q => n837);
   U834 : AO22X1 port map( IN1 => n5343, IN2 => RAMDIN1(23), IN3 => 
                           RAM_9_23_port, IN4 => n5337, Q => n838);
   U835 : AO22X1 port map( IN1 => n5344, IN2 => n2105, IN3 => RAM_9_24_port, 
                           IN4 => n5337, Q => n839);
   U836 : AO22X1 port map( IN1 => n5344, IN2 => RAMDIN1(25), IN3 => 
                           RAM_9_25_port, IN4 => n5337, Q => n840);
   U837 : AO22X1 port map( IN1 => n5344, IN2 => RAMDIN1(26), IN3 => 
                           RAM_9_26_port, IN4 => n5337, Q => n841);
   U838 : AO22X1 port map( IN1 => n5344, IN2 => RAMDIN1(27), IN3 => 
                           RAM_9_27_port, IN4 => n5337, Q => n842);
   U839 : AO22X1 port map( IN1 => RAMDIN1(28), IN2 => n5344, IN3 => 
                           RAM_9_28_port, IN4 => n5337, Q => n843);
   U840 : AO22X1 port map( IN1 => n5345, IN2 => RAMDIN1(29), IN3 => 
                           RAM_9_29_port, IN4 => n5337, Q => n844);
   U841 : AO22X1 port map( IN1 => n5345, IN2 => RAMDIN1(30), IN3 => 
                           RAM_9_30_port, IN4 => n5337, Q => n845);
   U842 : AO22X1 port map( IN1 => n5345, IN2 => RAMDIN1(31), IN3 => 
                           RAM_9_31_port, IN4 => n5337, Q => n846);
   U843 : AO22X1 port map( IN1 => n5345, IN2 => RAMDIN1(32), IN3 => 
                           RAM_9_32_port, IN4 => n5336, Q => n847);
   U844 : AO22X1 port map( IN1 => n5345, IN2 => RAMDIN1(33), IN3 => 
                           RAM_9_33_port, IN4 => n5336, Q => n848);
   U845 : AO22X1 port map( IN1 => n5346, IN2 => RAMDIN1(34), IN3 => 
                           RAM_9_34_port, IN4 => n5336, Q => n849);
   U846 : AO22X1 port map( IN1 => n5346, IN2 => RAMDIN1(35), IN3 => 
                           RAM_9_35_port, IN4 => n5336, Q => n850);
   U847 : AO22X1 port map( IN1 => n5346, IN2 => RAMDIN1(36), IN3 => 
                           RAM_9_36_port, IN4 => n5336, Q => n851);
   U848 : AO22X1 port map( IN1 => n5346, IN2 => n2558, IN3 => RAM_9_37_port, 
                           IN4 => n5336, Q => n852);
   U849 : AO22X1 port map( IN1 => n5346, IN2 => RAMDIN1(38), IN3 => 
                           RAM_9_38_port, IN4 => n5336, Q => n853);
   U850 : AO22X1 port map( IN1 => n5347, IN2 => RAMDIN1(39), IN3 => 
                           RAM_9_39_port, IN4 => n5336, Q => n854);
   U851 : AO22X1 port map( IN1 => n5347, IN2 => RAMDIN1(40), IN3 => 
                           RAM_9_40_port, IN4 => n5336, Q => n855);
   U852 : AO22X1 port map( IN1 => n5347, IN2 => n2507, IN3 => RAM_9_41_port, 
                           IN4 => n5336, Q => n856);
   U853 : AO22X1 port map( IN1 => n5347, IN2 => RAMDIN1(42), IN3 => 
                           RAM_9_42_port, IN4 => n5336, Q => n857);
   U854 : AO22X1 port map( IN1 => n5347, IN2 => n2560, IN3 => RAM_9_43_port, 
                           IN4 => n5336, Q => n858);
   U855 : AO22X1 port map( IN1 => RAMDIN1(44), IN2 => n5348, IN3 => 
                           RAM_9_44_port, IN4 => n5335, Q => n859);
   U856 : AO22X1 port map( IN1 => n5348, IN2 => RAMDIN1(45), IN3 => 
                           RAM_9_45_port, IN4 => n5335, Q => n860);
   U857 : AO22X1 port map( IN1 => RAMDIN1(46), IN2 => n5348, IN3 => 
                           RAM_9_46_port, IN4 => n5335, Q => n861);
   U858 : AO22X1 port map( IN1 => n5348, IN2 => RAMDIN1(47), IN3 => 
                           RAM_9_47_port, IN4 => n5335, Q => n862);
   U859 : AO22X1 port map( IN1 => n5348, IN2 => n2126, IN3 => RAM_9_48_port, 
                           IN4 => n5335, Q => n863);
   U860 : AO22X1 port map( IN1 => n5349, IN2 => RAMDIN1(49), IN3 => 
                           RAM_9_49_port, IN4 => n5335, Q => n864);
   U861 : AO22X1 port map( IN1 => n5349, IN2 => RAMDIN1(50), IN3 => 
                           RAM_9_50_port, IN4 => n5335, Q => n865);
   U862 : AO22X1 port map( IN1 => n5349, IN2 => RAMDIN1(51), IN3 => 
                           RAM_9_51_port, IN4 => n5335, Q => n866);
   U863 : AO22X1 port map( IN1 => n5349, IN2 => n2556, IN3 => RAM_9_52_port, 
                           IN4 => n5335, Q => n867);
   U864 : AO22X1 port map( IN1 => n5349, IN2 => RAMDIN1(53), IN3 => 
                           RAM_9_53_port, IN4 => n5335, Q => n868);
   U865 : AO22X1 port map( IN1 => n5350, IN2 => RAMDIN1(54), IN3 => 
                           RAM_9_54_port, IN4 => n5335, Q => n869);
   U866 : AO22X1 port map( IN1 => n5350, IN2 => RAMDIN1(55), IN3 => 
                           RAM_9_55_port, IN4 => n5335, Q => n870);
   U867 : AO22X1 port map( IN1 => n5350, IN2 => RAMDIN1(56), IN3 => 
                           RAM_9_56_port, IN4 => n5334, Q => n871);
   U868 : AO22X1 port map( IN1 => n5350, IN2 => RAMDIN1(57), IN3 => 
                           RAM_9_57_port, IN4 => n5334, Q => n872);
   U869 : AO22X1 port map( IN1 => n5350, IN2 => RAMDIN1(58), IN3 => 
                           RAM_9_58_port, IN4 => n5334, Q => n873);
   U870 : AO22X1 port map( IN1 => n5351, IN2 => RAMDIN1(59), IN3 => 
                           RAM_9_59_port, IN4 => n5334, Q => n874);
   U871 : AO22X1 port map( IN1 => n5351, IN2 => RAMDIN1(60), IN3 => 
                           RAM_9_60_port, IN4 => n5334, Q => n875);
   U872 : AO22X1 port map( IN1 => RAMDIN1(61), IN2 => n5351, IN3 => 
                           RAM_9_61_port, IN4 => n5334, Q => n876);
   U873 : AO22X1 port map( IN1 => n5351, IN2 => RAMDIN1(62), IN3 => 
                           RAM_9_62_port, IN4 => n5334, Q => n877);
   U874 : AO22X1 port map( IN1 => n5351, IN2 => RAMDIN1(63), IN3 => 
                           RAM_9_63_port, IN4 => n5334, Q => n878);
   U875 : AO22X1 port map( IN1 => n5352, IN2 => RAMDIN1(64), IN3 => 
                           RAM_9_64_port, IN4 => n5334, Q => n879);
   U876 : AO22X1 port map( IN1 => n5352, IN2 => RAMDIN1(65), IN3 => 
                           RAM_9_65_port, IN4 => n5334, Q => n880);
   U877 : AO22X1 port map( IN1 => n5352, IN2 => RAMDIN1(66), IN3 => 
                           RAM_9_66_port, IN4 => n5334, Q => n881);
   U878 : AO22X1 port map( IN1 => n5352, IN2 => RAMDIN1(67), IN3 => 
                           RAM_9_67_port, IN4 => n5334, Q => n882);
   U879 : AO22X1 port map( IN1 => n5352, IN2 => RAMDIN1(68), IN3 => 
                           RAM_9_68_port, IN4 => n5333, Q => n883);
   U880 : AO22X1 port map( IN1 => n5353, IN2 => RAMDIN1(69), IN3 => 
                           RAM_9_69_port, IN4 => n5333, Q => n884);
   U881 : AO22X1 port map( IN1 => n5353, IN2 => RAMDIN1(70), IN3 => 
                           RAM_9_70_port, IN4 => n5333, Q => n885);
   U882 : AO22X1 port map( IN1 => n5353, IN2 => RAMDIN1(71), IN3 => 
                           RAM_9_71_port, IN4 => n5333, Q => n886);
   U883 : AO22X1 port map( IN1 => n5353, IN2 => RAMDIN1(72), IN3 => 
                           RAM_9_72_port, IN4 => n5333, Q => n887);
   U884 : AO22X1 port map( IN1 => RAMDIN1(73), IN2 => n5353, IN3 => 
                           RAM_9_73_port, IN4 => n5333, Q => n888);
   U885 : AO22X1 port map( IN1 => n5354, IN2 => RAMDIN1(74), IN3 => 
                           RAM_9_74_port, IN4 => n5333, Q => n889);
   U886 : AO22X1 port map( IN1 => n5354, IN2 => RAMDIN1(75), IN3 => 
                           RAM_9_75_port, IN4 => n5333, Q => n890);
   U887 : AO22X1 port map( IN1 => n5354, IN2 => RAMDIN1(76), IN3 => 
                           RAM_9_76_port, IN4 => n5333, Q => n891);
   U888 : AO22X1 port map( IN1 => n5354, IN2 => RAMDIN1(77), IN3 => 
                           RAM_9_77_port, IN4 => n5333, Q => n892);
   U889 : AO22X1 port map( IN1 => n5354, IN2 => RAMDIN1(78), IN3 => 
                           RAM_9_78_port, IN4 => n5333, Q => n893);
   U890 : AO22X1 port map( IN1 => n5355, IN2 => RAMDIN1(79), IN3 => 
                           RAM_9_79_port, IN4 => n5333, Q => n894);
   U891 : AO22X1 port map( IN1 => RAMDIN1(80), IN2 => n5355, IN3 => 
                           RAM_9_80_port, IN4 => n5332, Q => n895);
   U892 : AO22X1 port map( IN1 => n5355, IN2 => RAMDIN1(81), IN3 => 
                           RAM_9_81_port, IN4 => n5332, Q => n896);
   U893 : AO22X1 port map( IN1 => n5355, IN2 => RAMDIN1(82), IN3 => 
                           RAM_9_82_port, IN4 => n5332, Q => n897);
   U894 : AO22X1 port map( IN1 => RAMDIN1(83), IN2 => n5355, IN3 => 
                           RAM_9_83_port, IN4 => n5332, Q => n898);
   U895 : AO22X1 port map( IN1 => RAMDIN1(84), IN2 => n5356, IN3 => 
                           RAM_9_84_port, IN4 => n5332, Q => n899);
   U896 : AO22X1 port map( IN1 => n5356, IN2 => RAMDIN1(85), IN3 => 
                           RAM_9_85_port, IN4 => n5332, Q => n900);
   U897 : AO22X1 port map( IN1 => n5356, IN2 => RAMDIN1(86), IN3 => 
                           RAM_9_86_port, IN4 => n5332, Q => n901);
   U898 : AO22X1 port map( IN1 => n5356, IN2 => RAMDIN1(87), IN3 => 
                           RAM_9_87_port, IN4 => n5332, Q => n902);
   U899 : AO22X1 port map( IN1 => RAMDIN1(88), IN2 => n5356, IN3 => 
                           RAM_9_88_port, IN4 => n5332, Q => n903);
   U900 : AO22X1 port map( IN1 => n5357, IN2 => RAMDIN1(89), IN3 => 
                           RAM_9_89_port, IN4 => n5332, Q => n904);
   U901 : AO22X1 port map( IN1 => n5357, IN2 => RAMDIN1(90), IN3 => 
                           RAM_9_90_port, IN4 => n5332, Q => n905);
   U902 : AO22X1 port map( IN1 => n5357, IN2 => RAMDIN1(91), IN3 => 
                           RAM_9_91_port, IN4 => n5332, Q => n906);
   U903 : AO22X1 port map( IN1 => n5357, IN2 => RAMDIN1(92), IN3 => 
                           RAM_9_92_port, IN4 => n5331, Q => n907);
   U904 : AO22X1 port map( IN1 => n5357, IN2 => RAMDIN1(93), IN3 => 
                           RAM_9_93_port, IN4 => n5331, Q => n908);
   U905 : AO22X1 port map( IN1 => n5358, IN2 => RAMDIN1(94), IN3 => 
                           RAM_9_94_port, IN4 => n5331, Q => n909);
   U906 : AO22X1 port map( IN1 => n5358, IN2 => RAMDIN1(95), IN3 => 
                           RAM_9_95_port, IN4 => n5331, Q => n910);
   U907 : AO22X1 port map( IN1 => n5358, IN2 => RAMDIN1(96), IN3 => 
                           RAM_9_96_port, IN4 => n5331, Q => n911);
   U908 : AO22X1 port map( IN1 => n5358, IN2 => RAMDIN1(97), IN3 => 
                           RAM_9_97_port, IN4 => n5331, Q => n912);
   U909 : AO22X1 port map( IN1 => n5358, IN2 => RAMDIN1(98), IN3 => 
                           RAM_9_98_port, IN4 => n5331, Q => n913);
   U910 : AO22X1 port map( IN1 => n5359, IN2 => n2102, IN3 => RAM_9_99_port, 
                           IN4 => n5331, Q => n914);
   U911 : AO22X1 port map( IN1 => n5359, IN2 => RAMDIN1(100), IN3 => 
                           RAM_9_100_port, IN4 => n5331, Q => n915);
   U912 : AO22X1 port map( IN1 => n5359, IN2 => RAMDIN1(101), IN3 => 
                           RAM_9_101_port, IN4 => n5331, Q => n916);
   U913 : AO22X1 port map( IN1 => n5359, IN2 => RAMDIN1(102), IN3 => 
                           RAM_9_102_port, IN4 => n5331, Q => n917);
   U914 : AO22X1 port map( IN1 => n5359, IN2 => RAMDIN1(103), IN3 => 
                           RAM_9_103_port, IN4 => n5331, Q => n918);
   U915 : AO22X1 port map( IN1 => n5360, IN2 => RAMDIN1(104), IN3 => 
                           RAM_9_104_port, IN4 => n5330, Q => n919);
   U916 : AO22X1 port map( IN1 => n5360, IN2 => RAMDIN1(105), IN3 => 
                           RAM_9_105_port, IN4 => n5330, Q => n920);
   U917 : AO22X1 port map( IN1 => n5360, IN2 => RAMDIN1(106), IN3 => 
                           RAM_9_106_port, IN4 => n5330, Q => n921);
   U918 : AO22X1 port map( IN1 => n5360, IN2 => RAMDIN1(107), IN3 => 
                           RAM_9_107_port, IN4 => n5330, Q => n922);
   U919 : AO22X1 port map( IN1 => n5360, IN2 => RAMDIN1(108), IN3 => 
                           RAM_9_108_port, IN4 => n5330, Q => n923);
   U920 : AO22X1 port map( IN1 => n5361, IN2 => RAMDIN1(109), IN3 => 
                           RAM_9_109_port, IN4 => n5330, Q => n924);
   U921 : AO22X1 port map( IN1 => RAMDIN1(110), IN2 => n5361, IN3 => 
                           RAM_9_110_port, IN4 => n5330, Q => n925);
   U922 : AO22X1 port map( IN1 => n5361, IN2 => RAMDIN1(111), IN3 => 
                           RAM_9_111_port, IN4 => n5330, Q => n926);
   U923 : AO22X1 port map( IN1 => RAMDIN1(112), IN2 => n5361, IN3 => 
                           RAM_9_112_port, IN4 => n5330, Q => n927);
   U924 : AO22X1 port map( IN1 => n5361, IN2 => RAMDIN1(113), IN3 => 
                           RAM_9_113_port, IN4 => n5330, Q => n928);
   U925 : AO22X1 port map( IN1 => n5362, IN2 => RAMDIN1(114), IN3 => 
                           RAM_9_114_port, IN4 => n5330, Q => n929);
   U926 : AO22X1 port map( IN1 => n5362, IN2 => RAMDIN1(115), IN3 => 
                           RAM_9_115_port, IN4 => n5330, Q => n930);
   U927 : AO22X1 port map( IN1 => n5362, IN2 => RAMDIN1(116), IN3 => 
                           RAM_9_116_port, IN4 => n5329, Q => n931);
   U928 : AO22X1 port map( IN1 => n5362, IN2 => RAMDIN1(117), IN3 => 
                           RAM_9_117_port, IN4 => n5329, Q => n932);
   U929 : AO22X1 port map( IN1 => n5362, IN2 => RAMDIN1(118), IN3 => 
                           RAM_9_118_port, IN4 => n5329, Q => n933);
   U930 : AO22X1 port map( IN1 => n5363, IN2 => RAMDIN1(119), IN3 => 
                           RAM_9_119_port, IN4 => n5329, Q => n934);
   U931 : AO22X1 port map( IN1 => n5363, IN2 => RAMDIN1(120), IN3 => 
                           RAM_9_120_port, IN4 => n5329, Q => n935);
   U932 : AO22X1 port map( IN1 => n5363, IN2 => RAMDIN1(121), IN3 => 
                           RAM_9_121_port, IN4 => n5329, Q => n936);
   U933 : AO22X1 port map( IN1 => n5363, IN2 => RAMDIN1(122), IN3 => 
                           RAM_9_122_port, IN4 => n5329, Q => n937);
   U934 : AO22X1 port map( IN1 => n5363, IN2 => RAMDIN1(123), IN3 => 
                           RAM_9_123_port, IN4 => n5329, Q => n938);
   U935 : AO22X1 port map( IN1 => n5364, IN2 => RAMDIN1(124), IN3 => 
                           RAM_9_124_port, IN4 => n5329, Q => n939);
   U936 : AO22X1 port map( IN1 => n5364, IN2 => RAMDIN1(125), IN3 => 
                           RAM_9_125_port, IN4 => n5329, Q => n940);
   U937 : AO22X1 port map( IN1 => n5364, IN2 => RAMDIN1(126), IN3 => 
                           RAM_9_126_port, IN4 => n5329, Q => n941);
   U938 : AO22X1 port map( IN1 => RAMDIN1(127), IN2 => n5364, IN3 => 
                           RAM_9_127_port, IN4 => n5329, Q => n942);
   U940 : AO22X1 port map( IN1 => n5301, IN2 => RAMDIN1(0), IN3 => RAM_8_0_port
                           , IN4 => n5297, Q => n943);
   U941 : AO22X1 port map( IN1 => n5300, IN2 => RAMDIN1(1), IN3 => RAM_8_1_port
                           , IN4 => n5297, Q => n944);
   U942 : AO22X1 port map( IN1 => n5298, IN2 => RAMDIN1(2), IN3 => RAM_8_2_port
                           , IN4 => n5297, Q => n945);
   U943 : AO22X1 port map( IN1 => n5298, IN2 => RAMDIN1(3), IN3 => RAM_8_3_port
                           , IN4 => n5297, Q => n946);
   U944 : AO22X1 port map( IN1 => n5320, IN2 => RAMDIN1(4), IN3 => RAM_8_4_port
                           , IN4 => n5297, Q => n947);
   U945 : AO22X1 port map( IN1 => n5322, IN2 => RAMDIN1(5), IN3 => RAM_8_5_port
                           , IN4 => n5297, Q => n948);
   U946 : AO22X1 port map( IN1 => n5321, IN2 => RAMDIN1(6), IN3 => RAM_8_6_port
                           , IN4 => n5297, Q => n949);
   U947 : AO22X1 port map( IN1 => n5320, IN2 => RAMDIN1(7), IN3 => RAM_8_7_port
                           , IN4 => n5297, Q => n950);
   U948 : AO22X1 port map( IN1 => n5322, IN2 => RAMDIN1(8), IN3 => RAM_8_8_port
                           , IN4 => n5296, Q => n951);
   U949 : AO22X1 port map( IN1 => n5322, IN2 => RAMDIN1(9), IN3 => RAM_8_9_port
                           , IN4 => n5296, Q => n952);
   U950 : AO22X1 port map( IN1 => n5321, IN2 => RAMDIN1(10), IN3 => 
                           RAM_8_10_port, IN4 => n5296, Q => n953);
   U951 : AO22X1 port map( IN1 => n5320, IN2 => RAMDIN1(11), IN3 => 
                           RAM_8_11_port, IN4 => n5296, Q => n954);
   U952 : AO22X1 port map( IN1 => n5322, IN2 => RAMDIN1(12), IN3 => 
                           RAM_8_12_port, IN4 => n5296, Q => n955);
   U953 : AO22X1 port map( IN1 => RAMDIN1(13), IN2 => n5321, IN3 => 
                           RAM_8_13_port, IN4 => n5296, Q => n956);
   U954 : AO22X1 port map( IN1 => RAMDIN1(14), IN2 => n5300, IN3 => 
                           RAM_8_14_port, IN4 => n5296, Q => n957);
   U955 : AO22X1 port map( IN1 => n5300, IN2 => RAMDIN1(15), IN3 => 
                           RAM_8_15_port, IN4 => n5296, Q => n958);
   U956 : AO22X1 port map( IN1 => RAMDIN1(16), IN2 => n5300, IN3 => 
                           RAM_8_16_port, IN4 => n5296, Q => n959);
   U957 : AO22X1 port map( IN1 => n5300, IN2 => RAMDIN1(17), IN3 => 
                           RAM_8_17_port, IN4 => n5296, Q => n960);
   U958 : AO22X1 port map( IN1 => n5300, IN2 => RAMDIN1(18), IN3 => 
                           RAM_8_18_port, IN4 => n5296, Q => n961);
   U959 : AO22X1 port map( IN1 => n5301, IN2 => RAMDIN1(19), IN3 => 
                           RAM_8_19_port, IN4 => n5296, Q => n962);
   U960 : AO22X1 port map( IN1 => n5301, IN2 => RAMDIN1(20), IN3 => 
                           RAM_8_20_port, IN4 => n5295, Q => n963);
   U961 : AO22X1 port map( IN1 => n5301, IN2 => RAMDIN1(21), IN3 => 
                           RAM_8_21_port, IN4 => n5295, Q => n964);
   U962 : AO22X1 port map( IN1 => n5301, IN2 => n2103, IN3 => RAM_8_22_port, 
                           IN4 => n5295, Q => n965);
   U963 : AO22X1 port map( IN1 => n5301, IN2 => RAMDIN1(23), IN3 => 
                           RAM_8_23_port, IN4 => n5295, Q => n966);
   U964 : AO22X1 port map( IN1 => n5302, IN2 => n2105, IN3 => RAM_8_24_port, 
                           IN4 => n5295, Q => n967);
   U965 : AO22X1 port map( IN1 => n5302, IN2 => RAMDIN1(25), IN3 => 
                           RAM_8_25_port, IN4 => n5295, Q => n968);
   U966 : AO22X1 port map( IN1 => n5302, IN2 => RAMDIN1(26), IN3 => 
                           RAM_8_26_port, IN4 => n5295, Q => n969);
   U967 : AO22X1 port map( IN1 => n5302, IN2 => RAMDIN1(27), IN3 => 
                           RAM_8_27_port, IN4 => n5295, Q => n970);
   U968 : AO22X1 port map( IN1 => RAMDIN1(28), IN2 => n5302, IN3 => 
                           RAM_8_28_port, IN4 => n5295, Q => n971);
   U969 : AO22X1 port map( IN1 => n5303, IN2 => RAMDIN1(29), IN3 => 
                           RAM_8_29_port, IN4 => n5295, Q => n972);
   U970 : AO22X1 port map( IN1 => n5303, IN2 => RAMDIN1(30), IN3 => 
                           RAM_8_30_port, IN4 => n5295, Q => n973);
   U971 : AO22X1 port map( IN1 => n5303, IN2 => RAMDIN1(31), IN3 => 
                           RAM_8_31_port, IN4 => n5295, Q => n974);
   U972 : AO22X1 port map( IN1 => n5303, IN2 => RAMDIN1(32), IN3 => 
                           RAM_8_32_port, IN4 => n5294, Q => n975);
   U973 : AO22X1 port map( IN1 => n5303, IN2 => RAMDIN1(33), IN3 => 
                           RAM_8_33_port, IN4 => n5294, Q => n976);
   U974 : AO22X1 port map( IN1 => n5304, IN2 => RAMDIN1(34), IN3 => 
                           RAM_8_34_port, IN4 => n5294, Q => n977);
   U975 : AO22X1 port map( IN1 => n5304, IN2 => RAMDIN1(35), IN3 => 
                           RAM_8_35_port, IN4 => n5294, Q => n978);
   U976 : AO22X1 port map( IN1 => n5304, IN2 => RAMDIN1(36), IN3 => 
                           RAM_8_36_port, IN4 => n5294, Q => n979);
   U977 : AO22X1 port map( IN1 => n5304, IN2 => n1, IN3 => RAM_8_37_port, IN4 
                           => n5294, Q => n980);
   U978 : AO22X1 port map( IN1 => n5304, IN2 => RAMDIN1(38), IN3 => 
                           RAM_8_38_port, IN4 => n5294, Q => n981);
   U979 : AO22X1 port map( IN1 => n5305, IN2 => RAMDIN1(39), IN3 => 
                           RAM_8_39_port, IN4 => n5294, Q => n982);
   U980 : AO22X1 port map( IN1 => n5305, IN2 => RAMDIN1(40), IN3 => 
                           RAM_8_40_port, IN4 => n5294, Q => n983);
   U981 : AO22X1 port map( IN1 => n5305, IN2 => n2507, IN3 => RAM_8_41_port, 
                           IN4 => n5294, Q => n984);
   U982 : AO22X1 port map( IN1 => n5305, IN2 => RAMDIN1(42), IN3 => 
                           RAM_8_42_port, IN4 => n5294, Q => n985);
   U983 : AO22X1 port map( IN1 => n5305, IN2 => n2101, IN3 => RAM_8_43_port, 
                           IN4 => n5294, Q => n986);
   U984 : AO22X1 port map( IN1 => RAMDIN1(44), IN2 => n5306, IN3 => 
                           RAM_8_44_port, IN4 => n5293, Q => n987);
   U985 : AO22X1 port map( IN1 => n5306, IN2 => RAMDIN1(45), IN3 => 
                           RAM_8_45_port, IN4 => n5293, Q => n988);
   U986 : AO22X1 port map( IN1 => RAMDIN1(46), IN2 => n5306, IN3 => 
                           RAM_8_46_port, IN4 => n5293, Q => n989);
   U987 : AO22X1 port map( IN1 => n5306, IN2 => RAMDIN1(47), IN3 => 
                           RAM_8_47_port, IN4 => n5293, Q => n990);
   U988 : AO22X1 port map( IN1 => n5306, IN2 => n2557, IN3 => RAM_8_48_port, 
                           IN4 => n5293, Q => n991);
   U989 : AO22X1 port map( IN1 => n5307, IN2 => RAMDIN1(49), IN3 => 
                           RAM_8_49_port, IN4 => n5293, Q => n992);
   U990 : AO22X1 port map( IN1 => n5307, IN2 => RAMDIN1(50), IN3 => 
                           RAM_8_50_port, IN4 => n5293, Q => n993);
   U991 : AO22X1 port map( IN1 => n5307, IN2 => RAMDIN1(51), IN3 => 
                           RAM_8_51_port, IN4 => n5293, Q => n994);
   U992 : AO22X1 port map( IN1 => n5307, IN2 => n2555, IN3 => RAM_8_52_port, 
                           IN4 => n5293, Q => n995);
   U993 : AO22X1 port map( IN1 => n5307, IN2 => RAMDIN1(53), IN3 => 
                           RAM_8_53_port, IN4 => n5293, Q => n996);
   U994 : AO22X1 port map( IN1 => n5308, IN2 => RAMDIN1(54), IN3 => 
                           RAM_8_54_port, IN4 => n5293, Q => n997);
   U995 : AO22X1 port map( IN1 => n5308, IN2 => RAMDIN1(55), IN3 => 
                           RAM_8_55_port, IN4 => n5293, Q => n998);
   U996 : AO22X1 port map( IN1 => n5308, IN2 => RAMDIN1(56), IN3 => 
                           RAM_8_56_port, IN4 => n5292, Q => n999);
   U997 : AO22X1 port map( IN1 => n5308, IN2 => RAMDIN1(57), IN3 => 
                           RAM_8_57_port, IN4 => n5292, Q => n1000);
   U998 : AO22X1 port map( IN1 => n5308, IN2 => RAMDIN1(58), IN3 => 
                           RAM_8_58_port, IN4 => n5292, Q => n1001);
   U999 : AO22X1 port map( IN1 => n5309, IN2 => RAMDIN1(59), IN3 => 
                           RAM_8_59_port, IN4 => n5292, Q => n1002);
   U1000 : AO22X1 port map( IN1 => n5309, IN2 => RAMDIN1(60), IN3 => 
                           RAM_8_60_port, IN4 => n5292, Q => n1003);
   U1001 : AO22X1 port map( IN1 => n5309, IN2 => RAMDIN1(61), IN3 => 
                           RAM_8_61_port, IN4 => n5292, Q => n1004);
   U1002 : AO22X1 port map( IN1 => n5309, IN2 => RAMDIN1(62), IN3 => 
                           RAM_8_62_port, IN4 => n5292, Q => n1005);
   U1003 : AO22X1 port map( IN1 => n5309, IN2 => RAMDIN1(63), IN3 => 
                           RAM_8_63_port, IN4 => n5292, Q => n1006);
   U1004 : AO22X1 port map( IN1 => n5310, IN2 => RAMDIN1(64), IN3 => 
                           RAM_8_64_port, IN4 => n5292, Q => n1007);
   U1005 : AO22X1 port map( IN1 => n5310, IN2 => RAMDIN1(65), IN3 => 
                           RAM_8_65_port, IN4 => n5292, Q => n1008);
   U1006 : AO22X1 port map( IN1 => n5310, IN2 => RAMDIN1(66), IN3 => 
                           RAM_8_66_port, IN4 => n5292, Q => n1009);
   U1007 : AO22X1 port map( IN1 => n5310, IN2 => RAMDIN1(67), IN3 => 
                           RAM_8_67_port, IN4 => n5292, Q => n1010);
   U1008 : AO22X1 port map( IN1 => n5310, IN2 => RAMDIN1(68), IN3 => 
                           RAM_8_68_port, IN4 => n5291, Q => n1011);
   U1009 : AO22X1 port map( IN1 => n5311, IN2 => RAMDIN1(69), IN3 => 
                           RAM_8_69_port, IN4 => n5291, Q => n1012);
   U1010 : AO22X1 port map( IN1 => n5311, IN2 => RAMDIN1(70), IN3 => 
                           RAM_8_70_port, IN4 => n5291, Q => n1013);
   U1011 : AO22X1 port map( IN1 => n5311, IN2 => RAMDIN1(71), IN3 => 
                           RAM_8_71_port, IN4 => n5291, Q => n1014);
   U1012 : AO22X1 port map( IN1 => n5311, IN2 => RAMDIN1(72), IN3 => 
                           RAM_8_72_port, IN4 => n5291, Q => n1015);
   U1013 : AO22X1 port map( IN1 => n5311, IN2 => RAMDIN1(73), IN3 => 
                           RAM_8_73_port, IN4 => n5291, Q => n1016);
   U1014 : AO22X1 port map( IN1 => n5312, IN2 => RAMDIN1(74), IN3 => 
                           RAM_8_74_port, IN4 => n5291, Q => n1017);
   U1015 : AO22X1 port map( IN1 => n5312, IN2 => RAMDIN1(75), IN3 => 
                           RAM_8_75_port, IN4 => n5291, Q => n1018);
   U1016 : AO22X1 port map( IN1 => n5312, IN2 => RAMDIN1(76), IN3 => 
                           RAM_8_76_port, IN4 => n5291, Q => n1019);
   U1017 : AO22X1 port map( IN1 => n5312, IN2 => RAMDIN1(77), IN3 => 
                           RAM_8_77_port, IN4 => n5291, Q => n1020);
   U1018 : AO22X1 port map( IN1 => n5312, IN2 => RAMDIN1(78), IN3 => 
                           RAM_8_78_port, IN4 => n5291, Q => n1021);
   U1019 : AO22X1 port map( IN1 => n5313, IN2 => RAMDIN1(79), IN3 => 
                           RAM_8_79_port, IN4 => n5291, Q => n1022);
   U1020 : AO22X1 port map( IN1 => RAMDIN1(80), IN2 => n5313, IN3 => 
                           RAM_8_80_port, IN4 => n5290, Q => n1023);
   U1021 : AO22X1 port map( IN1 => n5313, IN2 => RAMDIN1(81), IN3 => 
                           RAM_8_81_port, IN4 => n5290, Q => n1024);
   U1022 : AO22X1 port map( IN1 => n5313, IN2 => RAMDIN1(82), IN3 => 
                           RAM_8_82_port, IN4 => n5290, Q => n1025);
   U1023 : AO22X1 port map( IN1 => n5313, IN2 => RAMDIN1(83), IN3 => 
                           RAM_8_83_port, IN4 => n5290, Q => n1026);
   U1024 : AO22X1 port map( IN1 => n5314, IN2 => RAMDIN1(84), IN3 => 
                           RAM_8_84_port, IN4 => n5290, Q => n1027);
   U1025 : AO22X1 port map( IN1 => n5314, IN2 => RAMDIN1(85), IN3 => 
                           RAM_8_85_port, IN4 => n5290, Q => n1028);
   U1026 : AO22X1 port map( IN1 => n5314, IN2 => RAMDIN1(86), IN3 => 
                           RAM_8_86_port, IN4 => n5290, Q => n1029);
   U1027 : AO22X1 port map( IN1 => n5314, IN2 => RAMDIN1(87), IN3 => 
                           RAM_8_87_port, IN4 => n5290, Q => n1030);
   U1028 : AO22X1 port map( IN1 => RAMDIN1(88), IN2 => n5314, IN3 => 
                           RAM_8_88_port, IN4 => n5290, Q => n1031);
   U1029 : AO22X1 port map( IN1 => n5315, IN2 => RAMDIN1(89), IN3 => 
                           RAM_8_89_port, IN4 => n5290, Q => n1032);
   U1030 : AO22X1 port map( IN1 => n5315, IN2 => RAMDIN1(90), IN3 => 
                           RAM_8_90_port, IN4 => n5290, Q => n1033);
   U1031 : AO22X1 port map( IN1 => n5315, IN2 => RAMDIN1(91), IN3 => 
                           RAM_8_91_port, IN4 => n5290, Q => n1034);
   U1032 : AO22X1 port map( IN1 => n5315, IN2 => RAMDIN1(92), IN3 => 
                           RAM_8_92_port, IN4 => n5289, Q => n1035);
   U1033 : AO22X1 port map( IN1 => n5315, IN2 => RAMDIN1(93), IN3 => 
                           RAM_8_93_port, IN4 => n5289, Q => n1036);
   U1034 : AO22X1 port map( IN1 => n5316, IN2 => RAMDIN1(94), IN3 => 
                           RAM_8_94_port, IN4 => n5289, Q => n1037);
   U1035 : AO22X1 port map( IN1 => n5316, IN2 => RAMDIN1(95), IN3 => 
                           RAM_8_95_port, IN4 => n5289, Q => n1038);
   U1036 : AO22X1 port map( IN1 => n5316, IN2 => RAMDIN1(96), IN3 => 
                           RAM_8_96_port, IN4 => n5289, Q => n1039);
   U1037 : AO22X1 port map( IN1 => n5316, IN2 => RAMDIN1(97), IN3 => 
                           RAM_8_97_port, IN4 => n5289, Q => n1040);
   U1038 : AO22X1 port map( IN1 => n5316, IN2 => RAMDIN1(98), IN3 => 
                           RAM_8_98_port, IN4 => n5289, Q => n1041);
   U1039 : AO22X1 port map( IN1 => n5317, IN2 => n2502, IN3 => RAM_8_99_port, 
                           IN4 => n5289, Q => n1042);
   U1040 : AO22X1 port map( IN1 => n5317, IN2 => RAMDIN1(100), IN3 => 
                           RAM_8_100_port, IN4 => n5289, Q => n1043);
   U1041 : AO22X1 port map( IN1 => n5317, IN2 => RAMDIN1(101), IN3 => 
                           RAM_8_101_port, IN4 => n5289, Q => n1044);
   U1042 : AO22X1 port map( IN1 => n5317, IN2 => RAMDIN1(102), IN3 => 
                           RAM_8_102_port, IN4 => n5289, Q => n1045);
   U1043 : AO22X1 port map( IN1 => n5317, IN2 => RAMDIN1(103), IN3 => 
                           RAM_8_103_port, IN4 => n5289, Q => n1046);
   U1044 : AO22X1 port map( IN1 => n5318, IN2 => RAMDIN1(104), IN3 => 
                           RAM_8_104_port, IN4 => n5288, Q => n1047);
   U1045 : AO22X1 port map( IN1 => n5318, IN2 => RAMDIN1(105), IN3 => 
                           RAM_8_105_port, IN4 => n5288, Q => n1048);
   U1046 : AO22X1 port map( IN1 => n5318, IN2 => RAMDIN1(106), IN3 => 
                           RAM_8_106_port, IN4 => n5288, Q => n1049);
   U1047 : AO22X1 port map( IN1 => n5318, IN2 => RAMDIN1(107), IN3 => 
                           RAM_8_107_port, IN4 => n5288, Q => n1050);
   U1048 : AO22X1 port map( IN1 => n5318, IN2 => RAMDIN1(108), IN3 => 
                           RAM_8_108_port, IN4 => n5288, Q => n1051);
   U1049 : AO22X1 port map( IN1 => n5319, IN2 => RAMDIN1(109), IN3 => 
                           RAM_8_109_port, IN4 => n5288, Q => n1052);
   U1050 : AO22X1 port map( IN1 => RAMDIN1(110), IN2 => n5319, IN3 => 
                           RAM_8_110_port, IN4 => n5288, Q => n1053);
   U1051 : AO22X1 port map( IN1 => n5319, IN2 => RAMDIN1(111), IN3 => 
                           RAM_8_111_port, IN4 => n5288, Q => n1054);
   U1052 : AO22X1 port map( IN1 => RAMDIN1(112), IN2 => n5319, IN3 => 
                           RAM_8_112_port, IN4 => n5288, Q => n1055);
   U1053 : AO22X1 port map( IN1 => n5319, IN2 => RAMDIN1(113), IN3 => 
                           RAM_8_113_port, IN4 => n5288, Q => n1056);
   U1054 : AO22X1 port map( IN1 => n5320, IN2 => RAMDIN1(114), IN3 => 
                           RAM_8_114_port, IN4 => n5288, Q => n1057);
   U1055 : AO22X1 port map( IN1 => n5320, IN2 => RAMDIN1(115), IN3 => 
                           RAM_8_115_port, IN4 => n5288, Q => n1058);
   U1056 : AO22X1 port map( IN1 => n5320, IN2 => RAMDIN1(116), IN3 => 
                           RAM_8_116_port, IN4 => n5287, Q => n1059);
   U1057 : AO22X1 port map( IN1 => n5320, IN2 => RAMDIN1(117), IN3 => 
                           RAM_8_117_port, IN4 => n5287, Q => n1060);
   U1058 : AO22X1 port map( IN1 => n5320, IN2 => RAMDIN1(118), IN3 => 
                           RAM_8_118_port, IN4 => n5287, Q => n1061);
   U1059 : AO22X1 port map( IN1 => n5321, IN2 => RAMDIN1(119), IN3 => 
                           RAM_8_119_port, IN4 => n5287, Q => n1062);
   U1060 : AO22X1 port map( IN1 => n5321, IN2 => RAMDIN1(120), IN3 => 
                           RAM_8_120_port, IN4 => n5287, Q => n1063);
   U1061 : AO22X1 port map( IN1 => n5321, IN2 => RAMDIN1(121), IN3 => 
                           RAM_8_121_port, IN4 => n5287, Q => n1064);
   U1062 : AO22X1 port map( IN1 => n5321, IN2 => RAMDIN1(122), IN3 => 
                           RAM_8_122_port, IN4 => n5287, Q => n1065);
   U1063 : AO22X1 port map( IN1 => n5321, IN2 => RAMDIN1(123), IN3 => 
                           RAM_8_123_port, IN4 => n5287, Q => n1066);
   U1064 : AO22X1 port map( IN1 => n5322, IN2 => RAMDIN1(124), IN3 => 
                           RAM_8_124_port, IN4 => n5287, Q => n1067);
   U1065 : AO22X1 port map( IN1 => n5322, IN2 => RAMDIN1(125), IN3 => 
                           RAM_8_125_port, IN4 => n5287, Q => n1068);
   U1066 : AO22X1 port map( IN1 => n5322, IN2 => RAMDIN1(126), IN3 => 
                           RAM_8_126_port, IN4 => n5287, Q => n1069);
   U1067 : AO22X1 port map( IN1 => RAMDIN1(127), IN2 => n5322, IN3 => 
                           RAM_8_127_port, IN4 => n5287, Q => n1070);
   U1070 : AO22X1 port map( IN1 => n5259, IN2 => RAMDIN1(0), IN3 => 
                           RAM_7_0_port, IN4 => n5255, Q => n1071);
   U1071 : AO22X1 port map( IN1 => n5258, IN2 => RAMDIN1(1), IN3 => 
                           RAM_7_1_port, IN4 => n5255, Q => n1072);
   U1072 : AO22X1 port map( IN1 => n5256, IN2 => RAMDIN1(2), IN3 => 
                           RAM_7_2_port, IN4 => n5255, Q => n1073);
   U1073 : AO22X1 port map( IN1 => n5256, IN2 => RAMDIN1(3), IN3 => 
                           RAM_7_3_port, IN4 => n5255, Q => n1074);
   U1074 : AO22X1 port map( IN1 => n5278, IN2 => RAMDIN1(4), IN3 => 
                           RAM_7_4_port, IN4 => n5255, Q => n1075);
   U1075 : AO22X1 port map( IN1 => n5280, IN2 => RAMDIN1(5), IN3 => 
                           RAM_7_5_port, IN4 => n5255, Q => n1076);
   U1076 : AO22X1 port map( IN1 => n5279, IN2 => RAMDIN1(6), IN3 => 
                           RAM_7_6_port, IN4 => n5255, Q => n1077);
   U1077 : AO22X1 port map( IN1 => n5278, IN2 => RAMDIN1(7), IN3 => 
                           RAM_7_7_port, IN4 => n5255, Q => n1078);
   U1078 : AO22X1 port map( IN1 => n5280, IN2 => RAMDIN1(8), IN3 => 
                           RAM_7_8_port, IN4 => n5254, Q => n1079);
   U1079 : AO22X1 port map( IN1 => n5280, IN2 => RAMDIN1(9), IN3 => 
                           RAM_7_9_port, IN4 => n5254, Q => n1080);
   U1080 : AO22X1 port map( IN1 => n5279, IN2 => RAMDIN1(10), IN3 => 
                           RAM_7_10_port, IN4 => n5254, Q => n1081);
   U1081 : AO22X1 port map( IN1 => n5278, IN2 => RAMDIN1(11), IN3 => 
                           RAM_7_11_port, IN4 => n5254, Q => n1082);
   U1082 : AO22X1 port map( IN1 => n5280, IN2 => RAMDIN1(12), IN3 => 
                           RAM_7_12_port, IN4 => n5254, Q => n1083);
   U1083 : AO22X1 port map( IN1 => RAMDIN1(13), IN2 => n5279, IN3 => 
                           RAM_7_13_port, IN4 => n5254, Q => n1084);
   U1084 : AO22X1 port map( IN1 => RAMDIN1(14), IN2 => n5258, IN3 => 
                           RAM_7_14_port, IN4 => n5254, Q => n1085);
   U1085 : AO22X1 port map( IN1 => n5258, IN2 => RAMDIN1(15), IN3 => 
                           RAM_7_15_port, IN4 => n5254, Q => n1086);
   U1086 : AO22X1 port map( IN1 => RAMDIN1(16), IN2 => n5258, IN3 => 
                           RAM_7_16_port, IN4 => n5254, Q => n1087);
   U1087 : AO22X1 port map( IN1 => n5258, IN2 => RAMDIN1(17), IN3 => 
                           RAM_7_17_port, IN4 => n5254, Q => n1088);
   U1088 : AO22X1 port map( IN1 => n5258, IN2 => RAMDIN1(18), IN3 => 
                           RAM_7_18_port, IN4 => n5254, Q => n1089);
   U1089 : AO22X1 port map( IN1 => n5259, IN2 => RAMDIN1(19), IN3 => 
                           RAM_7_19_port, IN4 => n5254, Q => n1090);
   U1090 : AO22X1 port map( IN1 => n5259, IN2 => RAMDIN1(20), IN3 => 
                           RAM_7_20_port, IN4 => n5253, Q => n1091);
   U1091 : AO22X1 port map( IN1 => n5259, IN2 => RAMDIN1(21), IN3 => 
                           RAM_7_21_port, IN4 => n5253, Q => n1092);
   U1092 : AO22X1 port map( IN1 => n5259, IN2 => n2249, IN3 => RAM_7_22_port, 
                           IN4 => n5253, Q => n1093);
   U1093 : AO22X1 port map( IN1 => n5259, IN2 => RAMDIN1(23), IN3 => 
                           RAM_7_23_port, IN4 => n5253, Q => n1094);
   U1094 : AO22X1 port map( IN1 => n5260, IN2 => n2106, IN3 => RAM_7_24_port, 
                           IN4 => n5253, Q => n1095);
   U1095 : AO22X1 port map( IN1 => n5260, IN2 => RAMDIN1(25), IN3 => 
                           RAM_7_25_port, IN4 => n5253, Q => n1096);
   U1096 : AO22X1 port map( IN1 => n5260, IN2 => RAMDIN1(26), IN3 => 
                           RAM_7_26_port, IN4 => n5253, Q => n1097);
   U1097 : AO22X1 port map( IN1 => n5260, IN2 => RAMDIN1(27), IN3 => 
                           RAM_7_27_port, IN4 => n5253, Q => n1098);
   U1098 : AO22X1 port map( IN1 => RAMDIN1(28), IN2 => n5260, IN3 => 
                           RAM_7_28_port, IN4 => n5253, Q => n1099);
   U1099 : AO22X1 port map( IN1 => n5261, IN2 => RAMDIN1(29), IN3 => 
                           RAM_7_29_port, IN4 => n5253, Q => n1100);
   U1100 : AO22X1 port map( IN1 => n5261, IN2 => RAMDIN1(30), IN3 => 
                           RAM_7_30_port, IN4 => n5253, Q => n1101);
   U1101 : AO22X1 port map( IN1 => n5261, IN2 => RAMDIN1(31), IN3 => 
                           RAM_7_31_port, IN4 => n5253, Q => n1102);
   U1102 : AO22X1 port map( IN1 => n5261, IN2 => RAMDIN1(32), IN3 => 
                           RAM_7_32_port, IN4 => n5252, Q => n1103);
   U1103 : AO22X1 port map( IN1 => n5261, IN2 => RAMDIN1(33), IN3 => 
                           RAM_7_33_port, IN4 => n5252, Q => n1104);
   U1104 : AO22X1 port map( IN1 => n5262, IN2 => RAMDIN1(34), IN3 => 
                           RAM_7_34_port, IN4 => n5252, Q => n1105);
   U1105 : AO22X1 port map( IN1 => n5262, IN2 => RAMDIN1(35), IN3 => 
                           RAM_7_35_port, IN4 => n5252, Q => n1106);
   U1106 : AO22X1 port map( IN1 => n5262, IN2 => RAMDIN1(36), IN3 => 
                           RAM_7_36_port, IN4 => n5252, Q => n1107);
   U1107 : AO22X1 port map( IN1 => n5262, IN2 => n2558, IN3 => RAM_7_37_port, 
                           IN4 => n5252, Q => n1108);
   U1108 : AO22X1 port map( IN1 => n5262, IN2 => RAMDIN1(38), IN3 => 
                           RAM_7_38_port, IN4 => n5252, Q => n1109);
   U1109 : AO22X1 port map( IN1 => n5263, IN2 => RAMDIN1(39), IN3 => 
                           RAM_7_39_port, IN4 => n5252, Q => n1110);
   U1110 : AO22X1 port map( IN1 => n5263, IN2 => RAMDIN1(40), IN3 => 
                           RAM_7_40_port, IN4 => n5252, Q => n1111);
   U1111 : AO22X1 port map( IN1 => n5263, IN2 => n2506, IN3 => RAM_7_41_port, 
                           IN4 => n5252, Q => n1112);
   U1112 : AO22X1 port map( IN1 => n5263, IN2 => RAMDIN1(42), IN3 => 
                           RAM_7_42_port, IN4 => n5252, Q => n1113);
   U1113 : AO22X1 port map( IN1 => n5263, IN2 => n2101, IN3 => RAM_7_43_port, 
                           IN4 => n5252, Q => n1114);
   U1114 : AO22X1 port map( IN1 => RAMDIN1(44), IN2 => n5264, IN3 => 
                           RAM_7_44_port, IN4 => n5251, Q => n1115);
   U1115 : AO22X1 port map( IN1 => n5264, IN2 => RAMDIN1(45), IN3 => 
                           RAM_7_45_port, IN4 => n5251, Q => n1116);
   U1116 : AO22X1 port map( IN1 => RAMDIN1(46), IN2 => n5264, IN3 => 
                           RAM_7_46_port, IN4 => n5251, Q => n1117);
   U1117 : AO22X1 port map( IN1 => n5264, IN2 => RAMDIN1(47), IN3 => 
                           RAM_7_47_port, IN4 => n5251, Q => n1118);
   U1118 : AO22X1 port map( IN1 => n5264, IN2 => n2127, IN3 => RAM_7_48_port, 
                           IN4 => n5251, Q => n1119);
   U1119 : AO22X1 port map( IN1 => n5265, IN2 => RAMDIN1(49), IN3 => 
                           RAM_7_49_port, IN4 => n5251, Q => n1120);
   U1120 : AO22X1 port map( IN1 => n5265, IN2 => RAMDIN1(50), IN3 => 
                           RAM_7_50_port, IN4 => n5251, Q => n1121);
   U1121 : AO22X1 port map( IN1 => n5265, IN2 => RAMDIN1(51), IN3 => 
                           RAM_7_51_port, IN4 => n5251, Q => n1122);
   U1122 : AO22X1 port map( IN1 => n5265, IN2 => n2556, IN3 => RAM_7_52_port, 
                           IN4 => n5251, Q => n1123);
   U1123 : AO22X1 port map( IN1 => n5265, IN2 => RAMDIN1(53), IN3 => 
                           RAM_7_53_port, IN4 => n5251, Q => n1124);
   U1124 : AO22X1 port map( IN1 => n5266, IN2 => RAMDIN1(54), IN3 => 
                           RAM_7_54_port, IN4 => n5251, Q => n1125);
   U1125 : AO22X1 port map( IN1 => n5266, IN2 => RAMDIN1(55), IN3 => 
                           RAM_7_55_port, IN4 => n5251, Q => n1126);
   U1126 : AO22X1 port map( IN1 => n5266, IN2 => RAMDIN1(56), IN3 => 
                           RAM_7_56_port, IN4 => n5250, Q => n1127);
   U1127 : AO22X1 port map( IN1 => n5266, IN2 => RAMDIN1(57), IN3 => 
                           RAM_7_57_port, IN4 => n5250, Q => n1128);
   U1128 : AO22X1 port map( IN1 => n5266, IN2 => RAMDIN1(58), IN3 => 
                           RAM_7_58_port, IN4 => n5250, Q => n1129);
   U1129 : AO22X1 port map( IN1 => n5267, IN2 => RAMDIN1(59), IN3 => 
                           RAM_7_59_port, IN4 => n5250, Q => n1130);
   U1130 : AO22X1 port map( IN1 => n5267, IN2 => RAMDIN1(60), IN3 => 
                           RAM_7_60_port, IN4 => n5250, Q => n1131);
   U1131 : AO22X1 port map( IN1 => n5267, IN2 => RAMDIN1(61), IN3 => 
                           RAM_7_61_port, IN4 => n5250, Q => n1132);
   U1132 : AO22X1 port map( IN1 => n5267, IN2 => RAMDIN1(62), IN3 => 
                           RAM_7_62_port, IN4 => n5250, Q => n1133);
   U1133 : AO22X1 port map( IN1 => n5267, IN2 => RAMDIN1(63), IN3 => 
                           RAM_7_63_port, IN4 => n5250, Q => n1134);
   U1134 : AO22X1 port map( IN1 => n5268, IN2 => RAMDIN1(64), IN3 => 
                           RAM_7_64_port, IN4 => n5250, Q => n1135);
   U1135 : AO22X1 port map( IN1 => n5268, IN2 => RAMDIN1(65), IN3 => 
                           RAM_7_65_port, IN4 => n5250, Q => n1136);
   U1136 : AO22X1 port map( IN1 => n5268, IN2 => RAMDIN1(66), IN3 => 
                           RAM_7_66_port, IN4 => n5250, Q => n1137);
   U1137 : AO22X1 port map( IN1 => n5268, IN2 => RAMDIN1(67), IN3 => 
                           RAM_7_67_port, IN4 => n5250, Q => n1138);
   U1138 : AO22X1 port map( IN1 => n5268, IN2 => RAMDIN1(68), IN3 => 
                           RAM_7_68_port, IN4 => n5249, Q => n1139);
   U1139 : AO22X1 port map( IN1 => n5269, IN2 => RAMDIN1(69), IN3 => 
                           RAM_7_69_port, IN4 => n5249, Q => n1140);
   U1140 : AO22X1 port map( IN1 => n5269, IN2 => RAMDIN1(70), IN3 => 
                           RAM_7_70_port, IN4 => n5249, Q => n1141);
   U1141 : AO22X1 port map( IN1 => n5269, IN2 => RAMDIN1(71), IN3 => 
                           RAM_7_71_port, IN4 => n5249, Q => n1142);
   U1142 : AO22X1 port map( IN1 => n5269, IN2 => RAMDIN1(72), IN3 => 
                           RAM_7_72_port, IN4 => n5249, Q => n1143);
   U1143 : AO22X1 port map( IN1 => n5269, IN2 => RAMDIN1(73), IN3 => 
                           RAM_7_73_port, IN4 => n5249, Q => n1144);
   U1144 : AO22X1 port map( IN1 => n5270, IN2 => RAMDIN1(74), IN3 => 
                           RAM_7_74_port, IN4 => n5249, Q => n1145);
   U1145 : AO22X1 port map( IN1 => n5270, IN2 => RAMDIN1(75), IN3 => 
                           RAM_7_75_port, IN4 => n5249, Q => n1146);
   U1146 : AO22X1 port map( IN1 => n5270, IN2 => RAMDIN1(76), IN3 => 
                           RAM_7_76_port, IN4 => n5249, Q => n1147);
   U1147 : AO22X1 port map( IN1 => n5270, IN2 => RAMDIN1(77), IN3 => 
                           RAM_7_77_port, IN4 => n5249, Q => n1148);
   U1148 : AO22X1 port map( IN1 => n5270, IN2 => RAMDIN1(78), IN3 => 
                           RAM_7_78_port, IN4 => n5249, Q => n1149);
   U1149 : AO22X1 port map( IN1 => n5271, IN2 => RAMDIN1(79), IN3 => 
                           RAM_7_79_port, IN4 => n5249, Q => n1150);
   U1150 : AO22X1 port map( IN1 => RAMDIN1(80), IN2 => n5271, IN3 => 
                           RAM_7_80_port, IN4 => n5248, Q => n1151);
   U1151 : AO22X1 port map( IN1 => n5271, IN2 => RAMDIN1(81), IN3 => 
                           RAM_7_81_port, IN4 => n5248, Q => n1152);
   U1152 : AO22X1 port map( IN1 => n5271, IN2 => RAMDIN1(82), IN3 => 
                           RAM_7_82_port, IN4 => n5248, Q => n1153);
   U1153 : AO22X1 port map( IN1 => n5271, IN2 => RAMDIN1(83), IN3 => 
                           RAM_7_83_port, IN4 => n5248, Q => n1154);
   U1154 : AO22X1 port map( IN1 => n5272, IN2 => RAMDIN1(84), IN3 => 
                           RAM_7_84_port, IN4 => n5248, Q => n1155);
   U1155 : AO22X1 port map( IN1 => n5272, IN2 => RAMDIN1(85), IN3 => 
                           RAM_7_85_port, IN4 => n5248, Q => n1156);
   U1156 : AO22X1 port map( IN1 => n5272, IN2 => RAMDIN1(86), IN3 => 
                           RAM_7_86_port, IN4 => n5248, Q => n1157);
   U1157 : AO22X1 port map( IN1 => n5272, IN2 => RAMDIN1(87), IN3 => 
                           RAM_7_87_port, IN4 => n5248, Q => n1158);
   U1158 : AO22X1 port map( IN1 => RAMDIN1(88), IN2 => n5272, IN3 => 
                           RAM_7_88_port, IN4 => n5248, Q => n1159);
   U1159 : AO22X1 port map( IN1 => n5273, IN2 => RAMDIN1(89), IN3 => 
                           RAM_7_89_port, IN4 => n5248, Q => n1160);
   U1160 : AO22X1 port map( IN1 => n5273, IN2 => RAMDIN1(90), IN3 => 
                           RAM_7_90_port, IN4 => n5248, Q => n1161);
   U1161 : AO22X1 port map( IN1 => n5273, IN2 => RAMDIN1(91), IN3 => 
                           RAM_7_91_port, IN4 => n5248, Q => n1162);
   U1162 : AO22X1 port map( IN1 => n5273, IN2 => RAMDIN1(92), IN3 => 
                           RAM_7_92_port, IN4 => n5247, Q => n1163);
   U1163 : AO22X1 port map( IN1 => n5273, IN2 => RAMDIN1(93), IN3 => 
                           RAM_7_93_port, IN4 => n5247, Q => n1164);
   U1164 : AO22X1 port map( IN1 => n5274, IN2 => RAMDIN1(94), IN3 => 
                           RAM_7_94_port, IN4 => n5247, Q => n1165);
   U1165 : AO22X1 port map( IN1 => n5274, IN2 => RAMDIN1(95), IN3 => 
                           RAM_7_95_port, IN4 => n5247, Q => n1166);
   U1166 : AO22X1 port map( IN1 => n5274, IN2 => RAMDIN1(96), IN3 => 
                           RAM_7_96_port, IN4 => n5247, Q => n1167);
   U1167 : AO22X1 port map( IN1 => n5274, IN2 => RAMDIN1(97), IN3 => 
                           RAM_7_97_port, IN4 => n5247, Q => n1168);
   U1168 : AO22X1 port map( IN1 => n5274, IN2 => RAMDIN1(98), IN3 => 
                           RAM_7_98_port, IN4 => n5247, Q => n1169);
   U1169 : AO22X1 port map( IN1 => n5275, IN2 => n2503, IN3 => RAM_7_99_port, 
                           IN4 => n5247, Q => n1170);
   U1170 : AO22X1 port map( IN1 => n5275, IN2 => RAMDIN1(100), IN3 => 
                           RAM_7_100_port, IN4 => n5247, Q => n1171);
   U1171 : AO22X1 port map( IN1 => n5275, IN2 => RAMDIN1(101), IN3 => 
                           RAM_7_101_port, IN4 => n5247, Q => n1172);
   U1172 : AO22X1 port map( IN1 => n5275, IN2 => RAMDIN1(102), IN3 => 
                           RAM_7_102_port, IN4 => n5247, Q => n1173);
   U1173 : AO22X1 port map( IN1 => n5275, IN2 => RAMDIN1(103), IN3 => 
                           RAM_7_103_port, IN4 => n5247, Q => n1174);
   U1174 : AO22X1 port map( IN1 => n5276, IN2 => RAMDIN1(104), IN3 => 
                           RAM_7_104_port, IN4 => n5246, Q => n1175);
   U1175 : AO22X1 port map( IN1 => n5276, IN2 => RAMDIN1(105), IN3 => 
                           RAM_7_105_port, IN4 => n5246, Q => n1176);
   U1176 : AO22X1 port map( IN1 => n5276, IN2 => RAMDIN1(106), IN3 => 
                           RAM_7_106_port, IN4 => n5246, Q => n1177);
   U1177 : AO22X1 port map( IN1 => n5276, IN2 => RAMDIN1(107), IN3 => 
                           RAM_7_107_port, IN4 => n5246, Q => n1178);
   U1178 : AO22X1 port map( IN1 => n5276, IN2 => RAMDIN1(108), IN3 => 
                           RAM_7_108_port, IN4 => n5246, Q => n1179);
   U1179 : AO22X1 port map( IN1 => n5277, IN2 => RAMDIN1(109), IN3 => 
                           RAM_7_109_port, IN4 => n5246, Q => n1180);
   U1180 : AO22X1 port map( IN1 => RAMDIN1(110), IN2 => n5277, IN3 => 
                           RAM_7_110_port, IN4 => n5246, Q => n1181);
   U1181 : AO22X1 port map( IN1 => n5277, IN2 => RAMDIN1(111), IN3 => 
                           RAM_7_111_port, IN4 => n5246, Q => n1182);
   U1182 : AO22X1 port map( IN1 => RAMDIN1(112), IN2 => n5277, IN3 => 
                           RAM_7_112_port, IN4 => n5246, Q => n1183);
   U1183 : AO22X1 port map( IN1 => n5277, IN2 => RAMDIN1(113), IN3 => 
                           RAM_7_113_port, IN4 => n5246, Q => n1184);
   U1184 : AO22X1 port map( IN1 => n5278, IN2 => RAMDIN1(114), IN3 => 
                           RAM_7_114_port, IN4 => n5246, Q => n1185);
   U1185 : AO22X1 port map( IN1 => n5278, IN2 => RAMDIN1(115), IN3 => 
                           RAM_7_115_port, IN4 => n5246, Q => n1186);
   U1186 : AO22X1 port map( IN1 => n5278, IN2 => RAMDIN1(116), IN3 => 
                           RAM_7_116_port, IN4 => n5245, Q => n1187);
   U1187 : AO22X1 port map( IN1 => n5278, IN2 => RAMDIN1(117), IN3 => 
                           RAM_7_117_port, IN4 => n5245, Q => n1188);
   U1188 : AO22X1 port map( IN1 => n5278, IN2 => RAMDIN1(118), IN3 => 
                           RAM_7_118_port, IN4 => n5245, Q => n1189);
   U1189 : AO22X1 port map( IN1 => n5279, IN2 => RAMDIN1(119), IN3 => 
                           RAM_7_119_port, IN4 => n5245, Q => n1190);
   U1190 : AO22X1 port map( IN1 => n5279, IN2 => RAMDIN1(120), IN3 => 
                           RAM_7_120_port, IN4 => n5245, Q => n1191);
   U1191 : AO22X1 port map( IN1 => n5279, IN2 => RAMDIN1(121), IN3 => 
                           RAM_7_121_port, IN4 => n5245, Q => n1192);
   U1192 : AO22X1 port map( IN1 => n5279, IN2 => RAMDIN1(122), IN3 => 
                           RAM_7_122_port, IN4 => n5245, Q => n1193);
   U1193 : AO22X1 port map( IN1 => n5279, IN2 => RAMDIN1(123), IN3 => 
                           RAM_7_123_port, IN4 => n5245, Q => n1194);
   U1194 : AO22X1 port map( IN1 => n5280, IN2 => RAMDIN1(124), IN3 => 
                           RAM_7_124_port, IN4 => n5245, Q => n1195);
   U1195 : AO22X1 port map( IN1 => n5280, IN2 => RAMDIN1(125), IN3 => 
                           RAM_7_125_port, IN4 => n5245, Q => n1196);
   U1196 : AO22X1 port map( IN1 => n5280, IN2 => RAMDIN1(126), IN3 => 
                           RAM_7_126_port, IN4 => n5245, Q => n1197);
   U1197 : AO22X1 port map( IN1 => RAMDIN1(127), IN2 => n5280, IN3 => 
                           RAM_7_127_port, IN4 => n5245, Q => n1198);
   U1198 : AO22X1 port map( IN1 => n5217, IN2 => RAMDIN1(0), IN3 => 
                           RAM_6_0_port, IN4 => n5213, Q => n1199);
   U1199 : AO22X1 port map( IN1 => n5216, IN2 => RAMDIN1(1), IN3 => 
                           RAM_6_1_port, IN4 => n5213, Q => n1200);
   U1200 : AO22X1 port map( IN1 => n5214, IN2 => RAMDIN1(2), IN3 => 
                           RAM_6_2_port, IN4 => n5213, Q => n1201);
   U1201 : AO22X1 port map( IN1 => n5214, IN2 => RAMDIN1(3), IN3 => 
                           RAM_6_3_port, IN4 => n5213, Q => n1202);
   U1202 : AO22X1 port map( IN1 => n5236, IN2 => RAMDIN1(4), IN3 => 
                           RAM_6_4_port, IN4 => n5213, Q => n1203);
   U1203 : AO22X1 port map( IN1 => n5238, IN2 => RAMDIN1(5), IN3 => 
                           RAM_6_5_port, IN4 => n5213, Q => n1204);
   U1204 : AO22X1 port map( IN1 => n5237, IN2 => RAMDIN1(6), IN3 => 
                           RAM_6_6_port, IN4 => n5213, Q => n1205);
   U1205 : AO22X1 port map( IN1 => n5236, IN2 => RAMDIN1(7), IN3 => 
                           RAM_6_7_port, IN4 => n5213, Q => n1206);
   U1206 : AO22X1 port map( IN1 => n5238, IN2 => RAMDIN1(8), IN3 => 
                           RAM_6_8_port, IN4 => n5212, Q => n1207);
   U1207 : AO22X1 port map( IN1 => n5238, IN2 => RAMDIN1(9), IN3 => 
                           RAM_6_9_port, IN4 => n5212, Q => n1208);
   U1208 : AO22X1 port map( IN1 => n5237, IN2 => RAMDIN1(10), IN3 => 
                           RAM_6_10_port, IN4 => n5212, Q => n1209);
   U1209 : AO22X1 port map( IN1 => n5236, IN2 => RAMDIN1(11), IN3 => 
                           RAM_6_11_port, IN4 => n5212, Q => n1210);
   U1210 : AO22X1 port map( IN1 => n5238, IN2 => RAMDIN1(12), IN3 => 
                           RAM_6_12_port, IN4 => n5212, Q => n1211);
   U1211 : AO22X1 port map( IN1 => RAMDIN1(13), IN2 => n5237, IN3 => 
                           RAM_6_13_port, IN4 => n5212, Q => n1212);
   U1212 : AO22X1 port map( IN1 => RAMDIN1(14), IN2 => n5216, IN3 => 
                           RAM_6_14_port, IN4 => n5212, Q => n1213);
   U1213 : AO22X1 port map( IN1 => n5216, IN2 => RAMDIN1(15), IN3 => 
                           RAM_6_15_port, IN4 => n5212, Q => n1214);
   U1214 : AO22X1 port map( IN1 => RAMDIN1(16), IN2 => n5216, IN3 => 
                           RAM_6_16_port, IN4 => n5212, Q => n1215);
   U1215 : AO22X1 port map( IN1 => n5216, IN2 => RAMDIN1(17), IN3 => 
                           RAM_6_17_port, IN4 => n5212, Q => n1216);
   U1216 : AO22X1 port map( IN1 => n5216, IN2 => RAMDIN1(18), IN3 => 
                           RAM_6_18_port, IN4 => n5212, Q => n1217);
   U1217 : AO22X1 port map( IN1 => n5217, IN2 => RAMDIN1(19), IN3 => 
                           RAM_6_19_port, IN4 => n5212, Q => n1218);
   U1218 : AO22X1 port map( IN1 => n5217, IN2 => RAMDIN1(20), IN3 => 
                           RAM_6_20_port, IN4 => n5211, Q => n1219);
   U1219 : AO22X1 port map( IN1 => n5217, IN2 => RAMDIN1(21), IN3 => 
                           RAM_6_21_port, IN4 => n5211, Q => n1220);
   U1220 : AO22X1 port map( IN1 => n5217, IN2 => n2103, IN3 => RAM_6_22_port, 
                           IN4 => n5211, Q => n1221);
   U1221 : AO22X1 port map( IN1 => n5217, IN2 => RAMDIN1(23), IN3 => 
                           RAM_6_23_port, IN4 => n5211, Q => n1222);
   U1222 : AO22X1 port map( IN1 => n5218, IN2 => n2105, IN3 => RAM_6_24_port, 
                           IN4 => n5211, Q => n1223);
   U1223 : AO22X1 port map( IN1 => n5218, IN2 => RAMDIN1(25), IN3 => 
                           RAM_6_25_port, IN4 => n5211, Q => n1224);
   U1224 : AO22X1 port map( IN1 => n5218, IN2 => RAMDIN1(26), IN3 => 
                           RAM_6_26_port, IN4 => n5211, Q => n1225);
   U1225 : AO22X1 port map( IN1 => n5218, IN2 => RAMDIN1(27), IN3 => 
                           RAM_6_27_port, IN4 => n5211, Q => n1226);
   U1226 : AO22X1 port map( IN1 => RAMDIN1(28), IN2 => n5218, IN3 => 
                           RAM_6_28_port, IN4 => n5211, Q => n1227);
   U1227 : AO22X1 port map( IN1 => n5219, IN2 => RAMDIN1(29), IN3 => 
                           RAM_6_29_port, IN4 => n5211, Q => n1228);
   U1228 : AO22X1 port map( IN1 => n5219, IN2 => RAMDIN1(30), IN3 => 
                           RAM_6_30_port, IN4 => n5211, Q => n1229);
   U1229 : AO22X1 port map( IN1 => n5219, IN2 => RAMDIN1(31), IN3 => 
                           RAM_6_31_port, IN4 => n5211, Q => n1230);
   U1230 : AO22X1 port map( IN1 => n5219, IN2 => RAMDIN1(32), IN3 => 
                           RAM_6_32_port, IN4 => n5210, Q => n1231);
   U1231 : AO22X1 port map( IN1 => n5219, IN2 => RAMDIN1(33), IN3 => 
                           RAM_6_33_port, IN4 => n5210, Q => n1232);
   U1232 : AO22X1 port map( IN1 => n5220, IN2 => RAMDIN1(34), IN3 => 
                           RAM_6_34_port, IN4 => n5210, Q => n1233);
   U1233 : AO22X1 port map( IN1 => n5220, IN2 => RAMDIN1(35), IN3 => 
                           RAM_6_35_port, IN4 => n5210, Q => n1234);
   U1234 : AO22X1 port map( IN1 => n5220, IN2 => RAMDIN1(36), IN3 => 
                           RAM_6_36_port, IN4 => n5210, Q => n1235);
   U1235 : AO22X1 port map( IN1 => n5220, IN2 => n1, IN3 => RAM_6_37_port, IN4 
                           => n5210, Q => n1236);
   U1236 : AO22X1 port map( IN1 => n5220, IN2 => RAMDIN1(38), IN3 => 
                           RAM_6_38_port, IN4 => n5210, Q => n1237);
   U1237 : AO22X1 port map( IN1 => n5221, IN2 => RAMDIN1(39), IN3 => 
                           RAM_6_39_port, IN4 => n5210, Q => n1238);
   U1238 : AO22X1 port map( IN1 => n5221, IN2 => RAMDIN1(40), IN3 => 
                           RAM_6_40_port, IN4 => n5210, Q => n1239);
   U1239 : AO22X1 port map( IN1 => n5221, IN2 => n2104, IN3 => RAM_6_41_port, 
                           IN4 => n5210, Q => n1240);
   U1240 : AO22X1 port map( IN1 => n5221, IN2 => RAMDIN1(42), IN3 => 
                           RAM_6_42_port, IN4 => n5210, Q => n1241);
   U1241 : AO22X1 port map( IN1 => n5221, IN2 => n2101, IN3 => RAM_6_43_port, 
                           IN4 => n5210, Q => n1242);
   U1242 : AO22X1 port map( IN1 => RAMDIN1(44), IN2 => n5222, IN3 => 
                           RAM_6_44_port, IN4 => n5209, Q => n1243);
   U1243 : AO22X1 port map( IN1 => n5222, IN2 => RAMDIN1(45), IN3 => 
                           RAM_6_45_port, IN4 => n5209, Q => n1244);
   U1244 : AO22X1 port map( IN1 => RAMDIN1(46), IN2 => n5222, IN3 => 
                           RAM_6_46_port, IN4 => n5209, Q => n1245);
   U1245 : AO22X1 port map( IN1 => n5222, IN2 => RAMDIN1(47), IN3 => 
                           RAM_6_47_port, IN4 => n5209, Q => n1246);
   U1246 : AO22X1 port map( IN1 => n5222, IN2 => n2126, IN3 => RAM_6_48_port, 
                           IN4 => n5209, Q => n1247);
   U1247 : AO22X1 port map( IN1 => n5223, IN2 => RAMDIN1(49), IN3 => 
                           RAM_6_49_port, IN4 => n5209, Q => n1248);
   U1248 : AO22X1 port map( IN1 => n5223, IN2 => RAMDIN1(50), IN3 => 
                           RAM_6_50_port, IN4 => n5209, Q => n1249);
   U1249 : AO22X1 port map( IN1 => n5223, IN2 => RAMDIN1(51), IN3 => 
                           RAM_6_51_port, IN4 => n5209, Q => n1250);
   U1251 : AO22X1 port map( IN1 => n5223, IN2 => RAMDIN1(53), IN3 => 
                           RAM_6_53_port, IN4 => n5209, Q => n1252);
   U1252 : AO22X1 port map( IN1 => n5224, IN2 => RAMDIN1(54), IN3 => 
                           RAM_6_54_port, IN4 => n5209, Q => n1253);
   U1253 : AO22X1 port map( IN1 => n5224, IN2 => RAMDIN1(55), IN3 => 
                           RAM_6_55_port, IN4 => n5209, Q => n1254);
   U1254 : AO22X1 port map( IN1 => n5224, IN2 => RAMDIN1(56), IN3 => 
                           RAM_6_56_port, IN4 => n5208, Q => n1255);
   U1255 : AO22X1 port map( IN1 => n5224, IN2 => RAMDIN1(57), IN3 => 
                           RAM_6_57_port, IN4 => n5208, Q => n1256);
   U1256 : AO22X1 port map( IN1 => n5224, IN2 => RAMDIN1(58), IN3 => 
                           RAM_6_58_port, IN4 => n5208, Q => n1257);
   U1257 : AO22X1 port map( IN1 => n5225, IN2 => RAMDIN1(59), IN3 => 
                           RAM_6_59_port, IN4 => n5208, Q => n1258);
   U1258 : AO22X1 port map( IN1 => n5225, IN2 => RAMDIN1(60), IN3 => 
                           RAM_6_60_port, IN4 => n5208, Q => n1259);
   U1259 : AO22X1 port map( IN1 => n5225, IN2 => RAMDIN1(61), IN3 => 
                           RAM_6_61_port, IN4 => n5208, Q => n1260);
   U1260 : AO22X1 port map( IN1 => n5225, IN2 => RAMDIN1(62), IN3 => 
                           RAM_6_62_port, IN4 => n5208, Q => n1261);
   U1261 : AO22X1 port map( IN1 => n5225, IN2 => RAMDIN1(63), IN3 => 
                           RAM_6_63_port, IN4 => n5208, Q => n1262);
   U1262 : AO22X1 port map( IN1 => n5226, IN2 => RAMDIN1(64), IN3 => 
                           RAM_6_64_port, IN4 => n5208, Q => n1263);
   U1263 : AO22X1 port map( IN1 => n5226, IN2 => RAMDIN1(65), IN3 => 
                           RAM_6_65_port, IN4 => n5208, Q => n1264);
   U1264 : AO22X1 port map( IN1 => n5226, IN2 => RAMDIN1(66), IN3 => 
                           RAM_6_66_port, IN4 => n5208, Q => n1265);
   U1265 : AO22X1 port map( IN1 => n5226, IN2 => RAMDIN1(67), IN3 => 
                           RAM_6_67_port, IN4 => n5208, Q => n1266);
   U1266 : AO22X1 port map( IN1 => n5226, IN2 => RAMDIN1(68), IN3 => 
                           RAM_6_68_port, IN4 => n5207, Q => n1267);
   U1267 : AO22X1 port map( IN1 => n5227, IN2 => RAMDIN1(69), IN3 => 
                           RAM_6_69_port, IN4 => n5207, Q => n1268);
   U1268 : AO22X1 port map( IN1 => n5227, IN2 => RAMDIN1(70), IN3 => 
                           RAM_6_70_port, IN4 => n5207, Q => n1269);
   U1269 : AO22X1 port map( IN1 => n5227, IN2 => RAMDIN1(71), IN3 => 
                           RAM_6_71_port, IN4 => n5207, Q => n1270);
   U1270 : AO22X1 port map( IN1 => n5227, IN2 => RAMDIN1(72), IN3 => 
                           RAM_6_72_port, IN4 => n5207, Q => n1271);
   U1271 : AO22X1 port map( IN1 => n5227, IN2 => RAMDIN1(73), IN3 => 
                           RAM_6_73_port, IN4 => n5207, Q => n1272);
   U1272 : AO22X1 port map( IN1 => n5228, IN2 => RAMDIN1(74), IN3 => 
                           RAM_6_74_port, IN4 => n5207, Q => n1273);
   U1273 : AO22X1 port map( IN1 => n5228, IN2 => RAMDIN1(75), IN3 => 
                           RAM_6_75_port, IN4 => n5207, Q => n1274);
   U1274 : AO22X1 port map( IN1 => n5228, IN2 => RAMDIN1(76), IN3 => 
                           RAM_6_76_port, IN4 => n5207, Q => n1275);
   U1275 : AO22X1 port map( IN1 => n5228, IN2 => RAMDIN1(77), IN3 => 
                           RAM_6_77_port, IN4 => n5207, Q => n1276);
   U1276 : AO22X1 port map( IN1 => n5228, IN2 => RAMDIN1(78), IN3 => 
                           RAM_6_78_port, IN4 => n5207, Q => n1277);
   U1277 : AO22X1 port map( IN1 => n5229, IN2 => RAMDIN1(79), IN3 => 
                           RAM_6_79_port, IN4 => n5207, Q => n1278);
   U1278 : AO22X1 port map( IN1 => RAMDIN1(80), IN2 => n5229, IN3 => 
                           RAM_6_80_port, IN4 => n5206, Q => n1279);
   U1279 : AO22X1 port map( IN1 => n5229, IN2 => RAMDIN1(81), IN3 => 
                           RAM_6_81_port, IN4 => n5206, Q => n1280);
   U1280 : AO22X1 port map( IN1 => n5229, IN2 => RAMDIN1(82), IN3 => 
                           RAM_6_82_port, IN4 => n5206, Q => n1281);
   U1281 : AO22X1 port map( IN1 => n5229, IN2 => RAMDIN1(83), IN3 => 
                           RAM_6_83_port, IN4 => n5206, Q => n1282);
   U1282 : AO22X1 port map( IN1 => n5230, IN2 => RAMDIN1(84), IN3 => 
                           RAM_6_84_port, IN4 => n5206, Q => n1283);
   U1283 : AO22X1 port map( IN1 => n5230, IN2 => RAMDIN1(85), IN3 => 
                           RAM_6_85_port, IN4 => n5206, Q => n1284);
   U1284 : AO22X1 port map( IN1 => n5230, IN2 => RAMDIN1(86), IN3 => 
                           RAM_6_86_port, IN4 => n5206, Q => n1285);
   U1285 : AO22X1 port map( IN1 => n5230, IN2 => RAMDIN1(87), IN3 => 
                           RAM_6_87_port, IN4 => n5206, Q => n1286);
   U1286 : AO22X1 port map( IN1 => RAMDIN1(88), IN2 => n5230, IN3 => 
                           RAM_6_88_port, IN4 => n5206, Q => n1287);
   U1287 : AO22X1 port map( IN1 => n5231, IN2 => RAMDIN1(89), IN3 => 
                           RAM_6_89_port, IN4 => n5206, Q => n1288);
   U1288 : AO22X1 port map( IN1 => n5231, IN2 => RAMDIN1(90), IN3 => 
                           RAM_6_90_port, IN4 => n5206, Q => n1289);
   U1289 : AO22X1 port map( IN1 => n5231, IN2 => RAMDIN1(91), IN3 => 
                           RAM_6_91_port, IN4 => n5206, Q => n1290);
   U1290 : AO22X1 port map( IN1 => n5231, IN2 => RAMDIN1(92), IN3 => 
                           RAM_6_92_port, IN4 => n5205, Q => n1291);
   U1291 : AO22X1 port map( IN1 => n5231, IN2 => RAMDIN1(93), IN3 => 
                           RAM_6_93_port, IN4 => n5205, Q => n1292);
   U1292 : AO22X1 port map( IN1 => n5232, IN2 => RAMDIN1(94), IN3 => 
                           RAM_6_94_port, IN4 => n5205, Q => n1293);
   U1293 : AO22X1 port map( IN1 => n5232, IN2 => RAMDIN1(95), IN3 => 
                           RAM_6_95_port, IN4 => n5205, Q => n1294);
   U1294 : AO22X1 port map( IN1 => n5232, IN2 => RAMDIN1(96), IN3 => 
                           RAM_6_96_port, IN4 => n5205, Q => n1295);
   U1295 : AO22X1 port map( IN1 => n5232, IN2 => RAMDIN1(97), IN3 => 
                           RAM_6_97_port, IN4 => n5205, Q => n1296);
   U1296 : AO22X1 port map( IN1 => n5232, IN2 => RAMDIN1(98), IN3 => 
                           RAM_6_98_port, IN4 => n5205, Q => n1297);
   U1297 : AO22X1 port map( IN1 => n5233, IN2 => n2102, IN3 => RAM_6_99_port, 
                           IN4 => n5205, Q => n1298);
   U1298 : AO22X1 port map( IN1 => n5233, IN2 => RAMDIN1(100), IN3 => 
                           RAM_6_100_port, IN4 => n5205, Q => n1299);
   U1299 : AO22X1 port map( IN1 => n5233, IN2 => RAMDIN1(101), IN3 => 
                           RAM_6_101_port, IN4 => n5205, Q => n1300);
   U1300 : AO22X1 port map( IN1 => n5233, IN2 => RAMDIN1(102), IN3 => 
                           RAM_6_102_port, IN4 => n5205, Q => n1301);
   U1301 : AO22X1 port map( IN1 => n5233, IN2 => RAMDIN1(103), IN3 => 
                           RAM_6_103_port, IN4 => n5205, Q => n1302);
   U1302 : AO22X1 port map( IN1 => n5234, IN2 => RAMDIN1(104), IN3 => 
                           RAM_6_104_port, IN4 => n5204, Q => n1303);
   U1303 : AO22X1 port map( IN1 => n5234, IN2 => RAMDIN1(105), IN3 => 
                           RAM_6_105_port, IN4 => n5204, Q => n1304);
   U1304 : AO22X1 port map( IN1 => n5234, IN2 => RAMDIN1(106), IN3 => 
                           RAM_6_106_port, IN4 => n5204, Q => n1305);
   U1305 : AO22X1 port map( IN1 => n5234, IN2 => RAMDIN1(107), IN3 => 
                           RAM_6_107_port, IN4 => n5204, Q => n1306);
   U1306 : AO22X1 port map( IN1 => n5234, IN2 => RAMDIN1(108), IN3 => 
                           RAM_6_108_port, IN4 => n5204, Q => n1307);
   U1307 : AO22X1 port map( IN1 => n5235, IN2 => RAMDIN1(109), IN3 => 
                           RAM_6_109_port, IN4 => n5204, Q => n1308);
   U1308 : AO22X1 port map( IN1 => RAMDIN1(110), IN2 => n5235, IN3 => 
                           RAM_6_110_port, IN4 => n5204, Q => n1309);
   U1309 : AO22X1 port map( IN1 => n5235, IN2 => RAMDIN1(111), IN3 => 
                           RAM_6_111_port, IN4 => n5204, Q => n1310);
   U1310 : AO22X1 port map( IN1 => RAMDIN1(112), IN2 => n5235, IN3 => 
                           RAM_6_112_port, IN4 => n5204, Q => n1311);
   U1311 : AO22X1 port map( IN1 => n5235, IN2 => RAMDIN1(113), IN3 => 
                           RAM_6_113_port, IN4 => n5204, Q => n1312);
   U1312 : AO22X1 port map( IN1 => n5236, IN2 => RAMDIN1(114), IN3 => 
                           RAM_6_114_port, IN4 => n5204, Q => n1313);
   U1313 : AO22X1 port map( IN1 => n5236, IN2 => RAMDIN1(115), IN3 => 
                           RAM_6_115_port, IN4 => n5204, Q => n1314);
   U1314 : AO22X1 port map( IN1 => n5236, IN2 => RAMDIN1(116), IN3 => 
                           RAM_6_116_port, IN4 => n5203, Q => n1315);
   U1315 : AO22X1 port map( IN1 => n5236, IN2 => RAMDIN1(117), IN3 => 
                           RAM_6_117_port, IN4 => n5203, Q => n1316);
   U1316 : AO22X1 port map( IN1 => n5236, IN2 => RAMDIN1(118), IN3 => 
                           RAM_6_118_port, IN4 => n5203, Q => n1317);
   U1317 : AO22X1 port map( IN1 => n5237, IN2 => RAMDIN1(119), IN3 => 
                           RAM_6_119_port, IN4 => n5203, Q => n1318);
   U1318 : AO22X1 port map( IN1 => n5237, IN2 => RAMDIN1(120), IN3 => 
                           RAM_6_120_port, IN4 => n5203, Q => n1319);
   U1319 : AO22X1 port map( IN1 => n5237, IN2 => RAMDIN1(121), IN3 => 
                           RAM_6_121_port, IN4 => n5203, Q => n1320);
   U1320 : AO22X1 port map( IN1 => n5237, IN2 => RAMDIN1(122), IN3 => 
                           RAM_6_122_port, IN4 => n5203, Q => n1321);
   U1321 : AO22X1 port map( IN1 => n5237, IN2 => RAMDIN1(123), IN3 => 
                           RAM_6_123_port, IN4 => n5203, Q => n1322);
   U1322 : AO22X1 port map( IN1 => n5238, IN2 => RAMDIN1(124), IN3 => 
                           RAM_6_124_port, IN4 => n5203, Q => n1323);
   U1323 : AO22X1 port map( IN1 => n5238, IN2 => RAMDIN1(125), IN3 => 
                           RAM_6_125_port, IN4 => n5203, Q => n1324);
   U1324 : AO22X1 port map( IN1 => n5238, IN2 => RAMDIN1(126), IN3 => 
                           RAM_6_126_port, IN4 => n5203, Q => n1325);
   U1325 : AO22X1 port map( IN1 => RAMDIN1(127), IN2 => n5238, IN3 => 
                           RAM_6_127_port, IN4 => n5203, Q => n1326);
   U1326 : AO22X1 port map( IN1 => n5175, IN2 => RAMDIN1(0), IN3 => 
                           RAM_5_0_port, IN4 => n5171, Q => n1327);
   U1327 : AO22X1 port map( IN1 => n5174, IN2 => RAMDIN1(1), IN3 => 
                           RAM_5_1_port, IN4 => n5171, Q => n1328);
   U1328 : AO22X1 port map( IN1 => n5172, IN2 => RAMDIN1(2), IN3 => 
                           RAM_5_2_port, IN4 => n5171, Q => n1329);
   U1329 : AO22X1 port map( IN1 => n5172, IN2 => RAMDIN1(3), IN3 => 
                           RAM_5_3_port, IN4 => n5171, Q => n1330);
   U1330 : AO22X1 port map( IN1 => n5194, IN2 => RAMDIN1(4), IN3 => 
                           RAM_5_4_port, IN4 => n5171, Q => n1331);
   U1331 : AO22X1 port map( IN1 => n5196, IN2 => RAMDIN1(5), IN3 => 
                           RAM_5_5_port, IN4 => n5171, Q => n1332);
   U1332 : AO22X1 port map( IN1 => n5195, IN2 => RAMDIN1(6), IN3 => 
                           RAM_5_6_port, IN4 => n5171, Q => n1333);
   U1333 : AO22X1 port map( IN1 => n5194, IN2 => RAMDIN1(7), IN3 => 
                           RAM_5_7_port, IN4 => n5171, Q => n1334);
   U1334 : AO22X1 port map( IN1 => n5196, IN2 => RAMDIN1(8), IN3 => 
                           RAM_5_8_port, IN4 => n5170, Q => n1335);
   U1335 : AO22X1 port map( IN1 => n5196, IN2 => RAMDIN1(9), IN3 => 
                           RAM_5_9_port, IN4 => n5170, Q => n1336);
   U1336 : AO22X1 port map( IN1 => n5195, IN2 => RAMDIN1(10), IN3 => 
                           RAM_5_10_port, IN4 => n5170, Q => n1337);
   U1337 : AO22X1 port map( IN1 => n5194, IN2 => RAMDIN1(11), IN3 => 
                           RAM_5_11_port, IN4 => n5170, Q => n1338);
   U1338 : AO22X1 port map( IN1 => n5196, IN2 => RAMDIN1(12), IN3 => 
                           RAM_5_12_port, IN4 => n5170, Q => n1339);
   U1339 : AO22X1 port map( IN1 => RAMDIN1(13), IN2 => n5195, IN3 => 
                           RAM_5_13_port, IN4 => n5170, Q => n1340);
   U1340 : AO22X1 port map( IN1 => RAMDIN1(14), IN2 => n5174, IN3 => 
                           RAM_5_14_port, IN4 => n5170, Q => n1341);
   U1341 : AO22X1 port map( IN1 => n5174, IN2 => RAMDIN1(15), IN3 => 
                           RAM_5_15_port, IN4 => n5170, Q => n1342);
   U1342 : AO22X1 port map( IN1 => RAMDIN1(16), IN2 => n5174, IN3 => 
                           RAM_5_16_port, IN4 => n5170, Q => n1343);
   U1343 : AO22X1 port map( IN1 => n5174, IN2 => RAMDIN1(17), IN3 => 
                           RAM_5_17_port, IN4 => n5170, Q => n1344);
   U1344 : AO22X1 port map( IN1 => n5174, IN2 => RAMDIN1(18), IN3 => 
                           RAM_5_18_port, IN4 => n5170, Q => n1345);
   U1345 : AO22X1 port map( IN1 => n5175, IN2 => RAMDIN1(19), IN3 => 
                           RAM_5_19_port, IN4 => n5170, Q => n1346);
   U1346 : AO22X1 port map( IN1 => n5175, IN2 => RAMDIN1(20), IN3 => 
                           RAM_5_20_port, IN4 => n5169, Q => n1347);
   U1347 : AO22X1 port map( IN1 => n5175, IN2 => RAMDIN1(21), IN3 => 
                           RAM_5_21_port, IN4 => n5169, Q => n1348);
   U1348 : AO22X1 port map( IN1 => n5175, IN2 => n2248, IN3 => RAM_5_22_port, 
                           IN4 => n5169, Q => n1349);
   U1349 : AO22X1 port map( IN1 => n5175, IN2 => RAMDIN1(23), IN3 => 
                           RAM_5_23_port, IN4 => n5169, Q => n1350);
   U1350 : AO22X1 port map( IN1 => n5176, IN2 => n2200, IN3 => RAM_5_24_port, 
                           IN4 => n5169, Q => n1351);
   U1351 : AO22X1 port map( IN1 => n5176, IN2 => RAMDIN1(25), IN3 => 
                           RAM_5_25_port, IN4 => n5169, Q => n1352);
   U1352 : AO22X1 port map( IN1 => n5176, IN2 => RAMDIN1(26), IN3 => 
                           RAM_5_26_port, IN4 => n5169, Q => n1353);
   U1353 : AO22X1 port map( IN1 => n5176, IN2 => RAMDIN1(27), IN3 => 
                           RAM_5_27_port, IN4 => n5169, Q => n1354);
   U1354 : AO22X1 port map( IN1 => RAMDIN1(28), IN2 => n5176, IN3 => 
                           RAM_5_28_port, IN4 => n5169, Q => n1355);
   U1355 : AO22X1 port map( IN1 => n5177, IN2 => RAMDIN1(29), IN3 => 
                           RAM_5_29_port, IN4 => n5169, Q => n1356);
   U1356 : AO22X1 port map( IN1 => n5177, IN2 => RAMDIN1(30), IN3 => 
                           RAM_5_30_port, IN4 => n5169, Q => n1357);
   U1357 : AO22X1 port map( IN1 => n5177, IN2 => RAMDIN1(31), IN3 => 
                           RAM_5_31_port, IN4 => n5169, Q => n1358);
   U1358 : AO22X1 port map( IN1 => n5177, IN2 => RAMDIN1(32), IN3 => 
                           RAM_5_32_port, IN4 => n5168, Q => n1359);
   U1359 : AO22X1 port map( IN1 => n5177, IN2 => RAMDIN1(33), IN3 => 
                           RAM_5_33_port, IN4 => n5168, Q => n1360);
   U1360 : AO22X1 port map( IN1 => n5178, IN2 => RAMDIN1(34), IN3 => 
                           RAM_5_34_port, IN4 => n5168, Q => n1361);
   U1361 : AO22X1 port map( IN1 => n5178, IN2 => RAMDIN1(35), IN3 => 
                           RAM_5_35_port, IN4 => n5168, Q => n1362);
   U1362 : AO22X1 port map( IN1 => n5178, IN2 => RAMDIN1(36), IN3 => 
                           RAM_5_36_port, IN4 => n5168, Q => n1363);
   U1363 : AO22X1 port map( IN1 => n5178, IN2 => n2559, IN3 => RAM_5_37_port, 
                           IN4 => n5168, Q => n1364);
   U1364 : AO22X1 port map( IN1 => n5178, IN2 => RAMDIN1(38), IN3 => 
                           RAM_5_38_port, IN4 => n5168, Q => n1365);
   U1365 : AO22X1 port map( IN1 => n5179, IN2 => RAMDIN1(39), IN3 => 
                           RAM_5_39_port, IN4 => n5168, Q => n1366);
   U1366 : AO22X1 port map( IN1 => n5179, IN2 => RAMDIN1(40), IN3 => 
                           RAM_5_40_port, IN4 => n5168, Q => n1367);
   U1367 : AO22X1 port map( IN1 => n5179, IN2 => n2506, IN3 => RAM_5_41_port, 
                           IN4 => n5168, Q => n1368);
   U1368 : AO22X1 port map( IN1 => n5179, IN2 => RAMDIN1(42), IN3 => 
                           RAM_5_42_port, IN4 => n5168, Q => n1369);
   U1369 : AO22X1 port map( IN1 => n5179, IN2 => n2561, IN3 => RAM_5_43_port, 
                           IN4 => n5168, Q => n1370);
   U1370 : AO22X1 port map( IN1 => RAMDIN1(44), IN2 => n5180, IN3 => 
                           RAM_5_44_port, IN4 => n5167, Q => n1371);
   U1371 : AO22X1 port map( IN1 => n5180, IN2 => RAMDIN1(45), IN3 => 
                           RAM_5_45_port, IN4 => n5167, Q => n1372);
   U1372 : AO22X1 port map( IN1 => RAMDIN1(46), IN2 => n5180, IN3 => 
                           RAM_5_46_port, IN4 => n5167, Q => n1373);
   U1373 : AO22X1 port map( IN1 => n5180, IN2 => RAMDIN1(47), IN3 => 
                           RAM_5_47_port, IN4 => n5167, Q => n1374);
   U1374 : AO22X1 port map( IN1 => n5180, IN2 => n2557, IN3 => RAM_5_48_port, 
                           IN4 => n5167, Q => n1375);
   U1375 : AO22X1 port map( IN1 => n5181, IN2 => RAMDIN1(49), IN3 => 
                           RAM_5_49_port, IN4 => n5167, Q => n1376);
   U1376 : AO22X1 port map( IN1 => n5181, IN2 => RAMDIN1(50), IN3 => 
                           RAM_5_50_port, IN4 => n5167, Q => n1377);
   U1377 : AO22X1 port map( IN1 => n5181, IN2 => RAMDIN1(51), IN3 => 
                           RAM_5_51_port, IN4 => n5167, Q => n1378);
   U1378 : AO22X1 port map( IN1 => n5181, IN2 => n2, IN3 => RAM_5_52_port, IN4 
                           => n5167, Q => n1379);
   U1379 : AO22X1 port map( IN1 => n5181, IN2 => RAMDIN1(53), IN3 => 
                           RAM_5_53_port, IN4 => n5167, Q => n1380);
   U1380 : AO22X1 port map( IN1 => n5182, IN2 => RAMDIN1(54), IN3 => 
                           RAM_5_54_port, IN4 => n5167, Q => n1381);
   U1381 : AO22X1 port map( IN1 => n5182, IN2 => RAMDIN1(55), IN3 => 
                           RAM_5_55_port, IN4 => n5167, Q => n1382);
   U1382 : AO22X1 port map( IN1 => n5182, IN2 => RAMDIN1(56), IN3 => 
                           RAM_5_56_port, IN4 => n5166, Q => n1383);
   U1383 : AO22X1 port map( IN1 => n5182, IN2 => RAMDIN1(57), IN3 => 
                           RAM_5_57_port, IN4 => n5166, Q => n1384);
   U1384 : AO22X1 port map( IN1 => n5182, IN2 => RAMDIN1(58), IN3 => 
                           RAM_5_58_port, IN4 => n5166, Q => n1385);
   U1385 : AO22X1 port map( IN1 => n5183, IN2 => RAMDIN1(59), IN3 => 
                           RAM_5_59_port, IN4 => n5166, Q => n1386);
   U1386 : AO22X1 port map( IN1 => n5183, IN2 => RAMDIN1(60), IN3 => 
                           RAM_5_60_port, IN4 => n5166, Q => n1387);
   U1387 : AO22X1 port map( IN1 => n5183, IN2 => RAMDIN1(61), IN3 => 
                           RAM_5_61_port, IN4 => n5166, Q => n1388);
   U1388 : AO22X1 port map( IN1 => n5183, IN2 => RAMDIN1(62), IN3 => 
                           RAM_5_62_port, IN4 => n5166, Q => n1389);
   U1389 : AO22X1 port map( IN1 => n5183, IN2 => RAMDIN1(63), IN3 => 
                           RAM_5_63_port, IN4 => n5166, Q => n1390);
   U1390 : AO22X1 port map( IN1 => n5184, IN2 => RAMDIN1(64), IN3 => 
                           RAM_5_64_port, IN4 => n5166, Q => n1391);
   U1391 : AO22X1 port map( IN1 => n5184, IN2 => RAMDIN1(65), IN3 => 
                           RAM_5_65_port, IN4 => n5166, Q => n1392);
   U1392 : AO22X1 port map( IN1 => n5184, IN2 => RAMDIN1(66), IN3 => 
                           RAM_5_66_port, IN4 => n5166, Q => n1393);
   U1393 : AO22X1 port map( IN1 => n5184, IN2 => RAMDIN1(67), IN3 => 
                           RAM_5_67_port, IN4 => n5166, Q => n1394);
   U1394 : AO22X1 port map( IN1 => n5184, IN2 => RAMDIN1(68), IN3 => 
                           RAM_5_68_port, IN4 => n5165, Q => n1395);
   U1395 : AO22X1 port map( IN1 => n5185, IN2 => RAMDIN1(69), IN3 => 
                           RAM_5_69_port, IN4 => n5165, Q => n1396);
   U1396 : AO22X1 port map( IN1 => n5185, IN2 => RAMDIN1(70), IN3 => 
                           RAM_5_70_port, IN4 => n5165, Q => n1397);
   U1397 : AO22X1 port map( IN1 => n5185, IN2 => RAMDIN1(71), IN3 => 
                           RAM_5_71_port, IN4 => n5165, Q => n1398);
   U1398 : AO22X1 port map( IN1 => n5185, IN2 => RAMDIN1(72), IN3 => 
                           RAM_5_72_port, IN4 => n5165, Q => n1399);
   U1399 : AO22X1 port map( IN1 => n5185, IN2 => RAMDIN1(73), IN3 => 
                           RAM_5_73_port, IN4 => n5165, Q => n1400);
   U1400 : AO22X1 port map( IN1 => n5186, IN2 => RAMDIN1(74), IN3 => 
                           RAM_5_74_port, IN4 => n5165, Q => n1401);
   U1401 : AO22X1 port map( IN1 => n5186, IN2 => RAMDIN1(75), IN3 => 
                           RAM_5_75_port, IN4 => n5165, Q => n1402);
   U1402 : AO22X1 port map( IN1 => n5186, IN2 => RAMDIN1(76), IN3 => 
                           RAM_5_76_port, IN4 => n5165, Q => n1403);
   U1403 : AO22X1 port map( IN1 => n5186, IN2 => RAMDIN1(77), IN3 => 
                           RAM_5_77_port, IN4 => n5165, Q => n1404);
   U1404 : AO22X1 port map( IN1 => n5186, IN2 => RAMDIN1(78), IN3 => 
                           RAM_5_78_port, IN4 => n5165, Q => n1405);
   U1405 : AO22X1 port map( IN1 => n5187, IN2 => RAMDIN1(79), IN3 => 
                           RAM_5_79_port, IN4 => n5165, Q => n1406);
   U1406 : AO22X1 port map( IN1 => RAMDIN1(80), IN2 => n5187, IN3 => 
                           RAM_5_80_port, IN4 => n5164, Q => n1407);
   U1407 : AO22X1 port map( IN1 => n5187, IN2 => RAMDIN1(81), IN3 => 
                           RAM_5_81_port, IN4 => n5164, Q => n1408);
   U1408 : AO22X1 port map( IN1 => n5187, IN2 => RAMDIN1(82), IN3 => 
                           RAM_5_82_port, IN4 => n5164, Q => n1409);
   U1409 : AO22X1 port map( IN1 => n5187, IN2 => RAMDIN1(83), IN3 => 
                           RAM_5_83_port, IN4 => n5164, Q => n1410);
   U1410 : AO22X1 port map( IN1 => n5188, IN2 => RAMDIN1(84), IN3 => 
                           RAM_5_84_port, IN4 => n5164, Q => n1411);
   U1411 : AO22X1 port map( IN1 => n5188, IN2 => RAMDIN1(85), IN3 => 
                           RAM_5_85_port, IN4 => n5164, Q => n1412);
   U1412 : AO22X1 port map( IN1 => n5188, IN2 => RAMDIN1(86), IN3 => 
                           RAM_5_86_port, IN4 => n5164, Q => n1413);
   U1413 : AO22X1 port map( IN1 => n5188, IN2 => RAMDIN1(87), IN3 => 
                           RAM_5_87_port, IN4 => n5164, Q => n1414);
   U1414 : AO22X1 port map( IN1 => RAMDIN1(88), IN2 => n5188, IN3 => 
                           RAM_5_88_port, IN4 => n5164, Q => n1415);
   U1415 : AO22X1 port map( IN1 => n5189, IN2 => RAMDIN1(89), IN3 => 
                           RAM_5_89_port, IN4 => n5164, Q => n1416);
   U1416 : AO22X1 port map( IN1 => n5189, IN2 => RAMDIN1(90), IN3 => 
                           RAM_5_90_port, IN4 => n5164, Q => n1417);
   U1417 : AO22X1 port map( IN1 => n5189, IN2 => RAMDIN1(91), IN3 => 
                           RAM_5_91_port, IN4 => n5164, Q => n1418);
   U1418 : AO22X1 port map( IN1 => n5189, IN2 => RAMDIN1(92), IN3 => 
                           RAM_5_92_port, IN4 => n5163, Q => n1419);
   U1419 : AO22X1 port map( IN1 => n5189, IN2 => RAMDIN1(93), IN3 => 
                           RAM_5_93_port, IN4 => n5163, Q => n1420);
   U1420 : AO22X1 port map( IN1 => n5190, IN2 => RAMDIN1(94), IN3 => 
                           RAM_5_94_port, IN4 => n5163, Q => n1421);
   U1421 : AO22X1 port map( IN1 => n5190, IN2 => RAMDIN1(95), IN3 => 
                           RAM_5_95_port, IN4 => n5163, Q => n1422);
   U1422 : AO22X1 port map( IN1 => n5190, IN2 => RAMDIN1(96), IN3 => 
                           RAM_5_96_port, IN4 => n5163, Q => n1423);
   U1423 : AO22X1 port map( IN1 => n5190, IN2 => RAMDIN1(97), IN3 => 
                           RAM_5_97_port, IN4 => n5163, Q => n1424);
   U1424 : AO22X1 port map( IN1 => n5190, IN2 => RAMDIN1(98), IN3 => 
                           RAM_5_98_port, IN4 => n5163, Q => n1425);
   U1425 : AO22X1 port map( IN1 => n5191, IN2 => n2502, IN3 => RAM_5_99_port, 
                           IN4 => n5163, Q => n1426);
   U1426 : AO22X1 port map( IN1 => n5191, IN2 => RAMDIN1(100), IN3 => 
                           RAM_5_100_port, IN4 => n5163, Q => n1427);
   U1427 : AO22X1 port map( IN1 => n5191, IN2 => RAMDIN1(101), IN3 => 
                           RAM_5_101_port, IN4 => n5163, Q => n1428);
   U1428 : AO22X1 port map( IN1 => n5191, IN2 => RAMDIN1(102), IN3 => 
                           RAM_5_102_port, IN4 => n5163, Q => n1429);
   U1429 : AO22X1 port map( IN1 => n5191, IN2 => RAMDIN1(103), IN3 => 
                           RAM_5_103_port, IN4 => n5163, Q => n1430);
   U1430 : AO22X1 port map( IN1 => n5192, IN2 => RAMDIN1(104), IN3 => 
                           RAM_5_104_port, IN4 => n5162, Q => n1431);
   U1431 : AO22X1 port map( IN1 => n5192, IN2 => RAMDIN1(105), IN3 => 
                           RAM_5_105_port, IN4 => n5162, Q => n1432);
   U1432 : AO22X1 port map( IN1 => n5192, IN2 => RAMDIN1(106), IN3 => 
                           RAM_5_106_port, IN4 => n5162, Q => n1433);
   U1433 : AO22X1 port map( IN1 => n5192, IN2 => RAMDIN1(107), IN3 => 
                           RAM_5_107_port, IN4 => n5162, Q => n1434);
   U1434 : AO22X1 port map( IN1 => n5192, IN2 => RAMDIN1(108), IN3 => 
                           RAM_5_108_port, IN4 => n5162, Q => n1435);
   U1435 : AO22X1 port map( IN1 => n5193, IN2 => RAMDIN1(109), IN3 => 
                           RAM_5_109_port, IN4 => n5162, Q => n1436);
   U1436 : AO22X1 port map( IN1 => RAMDIN1(110), IN2 => n5193, IN3 => 
                           RAM_5_110_port, IN4 => n5162, Q => n1437);
   U1437 : AO22X1 port map( IN1 => n5193, IN2 => RAMDIN1(111), IN3 => 
                           RAM_5_111_port, IN4 => n5162, Q => n1438);
   U1438 : AO22X1 port map( IN1 => RAMDIN1(112), IN2 => n5193, IN3 => 
                           RAM_5_112_port, IN4 => n5162, Q => n1439);
   U1439 : AO22X1 port map( IN1 => n5193, IN2 => RAMDIN1(113), IN3 => 
                           RAM_5_113_port, IN4 => n5162, Q => n1440);
   U1440 : AO22X1 port map( IN1 => n5194, IN2 => RAMDIN1(114), IN3 => 
                           RAM_5_114_port, IN4 => n5162, Q => n1441);
   U1441 : AO22X1 port map( IN1 => n5194, IN2 => RAMDIN1(115), IN3 => 
                           RAM_5_115_port, IN4 => n5162, Q => n1442);
   U1442 : AO22X1 port map( IN1 => n5194, IN2 => RAMDIN1(116), IN3 => 
                           RAM_5_116_port, IN4 => n5161, Q => n1443);
   U1443 : AO22X1 port map( IN1 => n5194, IN2 => RAMDIN1(117), IN3 => 
                           RAM_5_117_port, IN4 => n5161, Q => n1444);
   U1444 : AO22X1 port map( IN1 => n5194, IN2 => RAMDIN1(118), IN3 => 
                           RAM_5_118_port, IN4 => n5161, Q => n1445);
   U1445 : AO22X1 port map( IN1 => n5195, IN2 => RAMDIN1(119), IN3 => 
                           RAM_5_119_port, IN4 => n5161, Q => n1446);
   U1446 : AO22X1 port map( IN1 => n5195, IN2 => RAMDIN1(120), IN3 => 
                           RAM_5_120_port, IN4 => n5161, Q => n1447);
   U1447 : AO22X1 port map( IN1 => n5195, IN2 => RAMDIN1(121), IN3 => 
                           RAM_5_121_port, IN4 => n5161, Q => n1448);
   U1448 : AO22X1 port map( IN1 => n5195, IN2 => RAMDIN1(122), IN3 => 
                           RAM_5_122_port, IN4 => n5161, Q => n1449);
   U1449 : AO22X1 port map( IN1 => n5195, IN2 => RAMDIN1(123), IN3 => 
                           RAM_5_123_port, IN4 => n5161, Q => n1450);
   U1450 : AO22X1 port map( IN1 => n5196, IN2 => RAMDIN1(124), IN3 => 
                           RAM_5_124_port, IN4 => n5161, Q => n1451);
   U1451 : AO22X1 port map( IN1 => n5196, IN2 => RAMDIN1(125), IN3 => 
                           RAM_5_125_port, IN4 => n5161, Q => n1452);
   U1452 : AO22X1 port map( IN1 => n5196, IN2 => RAMDIN1(126), IN3 => 
                           RAM_5_126_port, IN4 => n5161, Q => n1453);
   U1453 : AO22X1 port map( IN1 => RAMDIN1(127), IN2 => n5196, IN3 => 
                           RAM_5_127_port, IN4 => n5161, Q => n1454);
   U1454 : AO22X1 port map( IN1 => n5133, IN2 => RAMDIN1(0), IN3 => 
                           RAM_4_0_port, IN4 => n5129, Q => n1455);
   U1455 : AO22X1 port map( IN1 => n5132, IN2 => RAMDIN1(1), IN3 => 
                           RAM_4_1_port, IN4 => n5129, Q => n1456);
   U1456 : AO22X1 port map( IN1 => n5130, IN2 => RAMDIN1(2), IN3 => 
                           RAM_4_2_port, IN4 => n5129, Q => n1457);
   U1457 : AO22X1 port map( IN1 => n5130, IN2 => RAMDIN1(3), IN3 => 
                           RAM_4_3_port, IN4 => n5129, Q => n1458);
   U1458 : AO22X1 port map( IN1 => n5152, IN2 => RAMDIN1(4), IN3 => 
                           RAM_4_4_port, IN4 => n5129, Q => n1459);
   U1459 : AO22X1 port map( IN1 => n5154, IN2 => RAMDIN1(5), IN3 => 
                           RAM_4_5_port, IN4 => n5129, Q => n1460);
   U1460 : AO22X1 port map( IN1 => n5153, IN2 => RAMDIN1(6), IN3 => 
                           RAM_4_6_port, IN4 => n5129, Q => n1461);
   U1461 : AO22X1 port map( IN1 => n5152, IN2 => RAMDIN1(7), IN3 => 
                           RAM_4_7_port, IN4 => n5129, Q => n1462);
   U1462 : AO22X1 port map( IN1 => n5154, IN2 => RAMDIN1(8), IN3 => 
                           RAM_4_8_port, IN4 => n5128, Q => n1463);
   U1463 : AO22X1 port map( IN1 => n5154, IN2 => RAMDIN1(9), IN3 => 
                           RAM_4_9_port, IN4 => n5128, Q => n1464);
   U1464 : AO22X1 port map( IN1 => n5153, IN2 => RAMDIN1(10), IN3 => 
                           RAM_4_10_port, IN4 => n5128, Q => n1465);
   U1465 : AO22X1 port map( IN1 => n5152, IN2 => RAMDIN1(11), IN3 => 
                           RAM_4_11_port, IN4 => n5128, Q => n1466);
   U1466 : AO22X1 port map( IN1 => n5154, IN2 => RAMDIN1(12), IN3 => 
                           RAM_4_12_port, IN4 => n5128, Q => n1467);
   U1467 : AO22X1 port map( IN1 => RAMDIN1(13), IN2 => n5153, IN3 => 
                           RAM_4_13_port, IN4 => n5128, Q => n1468);
   U1468 : AO22X1 port map( IN1 => RAMDIN1(14), IN2 => n5132, IN3 => 
                           RAM_4_14_port, IN4 => n5128, Q => n1469);
   U1469 : AO22X1 port map( IN1 => n5132, IN2 => RAMDIN1(15), IN3 => 
                           RAM_4_15_port, IN4 => n5128, Q => n1470);
   U1470 : AO22X1 port map( IN1 => RAMDIN1(16), IN2 => n5132, IN3 => 
                           RAM_4_16_port, IN4 => n5128, Q => n1471);
   U1471 : AO22X1 port map( IN1 => n5132, IN2 => RAMDIN1(17), IN3 => 
                           RAM_4_17_port, IN4 => n5128, Q => n1472);
   U1472 : AO22X1 port map( IN1 => n5132, IN2 => RAMDIN1(18), IN3 => 
                           RAM_4_18_port, IN4 => n5128, Q => n1473);
   U1473 : AO22X1 port map( IN1 => n5133, IN2 => RAMDIN1(19), IN3 => 
                           RAM_4_19_port, IN4 => n5128, Q => n1474);
   U1474 : AO22X1 port map( IN1 => n5133, IN2 => RAMDIN1(20), IN3 => 
                           RAM_4_20_port, IN4 => n5127, Q => n1475);
   U1475 : AO22X1 port map( IN1 => n5133, IN2 => RAMDIN1(21), IN3 => 
                           RAM_4_21_port, IN4 => n5127, Q => n1476);
   U1476 : AO22X1 port map( IN1 => n5133, IN2 => n2249, IN3 => RAM_4_22_port, 
                           IN4 => n5127, Q => n1477);
   U1477 : AO22X1 port map( IN1 => n5133, IN2 => RAMDIN1(23), IN3 => 
                           RAM_4_23_port, IN4 => n5127, Q => n1478);
   U1478 : AO22X1 port map( IN1 => n5134, IN2 => n2106, IN3 => RAM_4_24_port, 
                           IN4 => n5127, Q => n1479);
   U1479 : AO22X1 port map( IN1 => n5134, IN2 => RAMDIN1(25), IN3 => 
                           RAM_4_25_port, IN4 => n5127, Q => n1480);
   U1480 : AO22X1 port map( IN1 => n5134, IN2 => RAMDIN1(26), IN3 => 
                           RAM_4_26_port, IN4 => n5127, Q => n1481);
   U1481 : AO22X1 port map( IN1 => n5134, IN2 => RAMDIN1(27), IN3 => 
                           RAM_4_27_port, IN4 => n5127, Q => n1482);
   U1482 : AO22X1 port map( IN1 => RAMDIN1(28), IN2 => n5134, IN3 => 
                           RAM_4_28_port, IN4 => n5127, Q => n1483);
   U1483 : AO22X1 port map( IN1 => n5135, IN2 => RAMDIN1(29), IN3 => 
                           RAM_4_29_port, IN4 => n5127, Q => n1484);
   U1484 : AO22X1 port map( IN1 => n5135, IN2 => RAMDIN1(30), IN3 => 
                           RAM_4_30_port, IN4 => n5127, Q => n1485);
   U1485 : AO22X1 port map( IN1 => n5135, IN2 => RAMDIN1(31), IN3 => 
                           RAM_4_31_port, IN4 => n5127, Q => n1486);
   U1486 : AO22X1 port map( IN1 => n5135, IN2 => RAMDIN1(32), IN3 => 
                           RAM_4_32_port, IN4 => n5126, Q => n1487);
   U1487 : AO22X1 port map( IN1 => n5135, IN2 => RAMDIN1(33), IN3 => 
                           RAM_4_33_port, IN4 => n5126, Q => n1488);
   U1488 : AO22X1 port map( IN1 => n5136, IN2 => RAMDIN1(34), IN3 => 
                           RAM_4_34_port, IN4 => n5126, Q => n1489);
   U1489 : AO22X1 port map( IN1 => n5136, IN2 => RAMDIN1(35), IN3 => 
                           RAM_4_35_port, IN4 => n5126, Q => n1490);
   U1490 : AO22X1 port map( IN1 => n5136, IN2 => RAMDIN1(36), IN3 => 
                           RAM_4_36_port, IN4 => n5126, Q => n1491);
   U1491 : AO22X1 port map( IN1 => n5136, IN2 => n2558, IN3 => RAM_4_37_port, 
                           IN4 => n5126, Q => n1492);
   U1492 : AO22X1 port map( IN1 => n5136, IN2 => RAMDIN1(38), IN3 => 
                           RAM_4_38_port, IN4 => n5126, Q => n1493);
   U1493 : AO22X1 port map( IN1 => n5137, IN2 => RAMDIN1(39), IN3 => 
                           RAM_4_39_port, IN4 => n5126, Q => n1494);
   U1494 : AO22X1 port map( IN1 => n5137, IN2 => RAMDIN1(40), IN3 => 
                           RAM_4_40_port, IN4 => n5126, Q => n1495);
   U1495 : AO22X1 port map( IN1 => n5137, IN2 => n2104, IN3 => RAM_4_41_port, 
                           IN4 => n5126, Q => n1496);
   U1496 : AO22X1 port map( IN1 => n5137, IN2 => RAMDIN1(42), IN3 => 
                           RAM_4_42_port, IN4 => n5126, Q => n1497);
   U1497 : AO22X1 port map( IN1 => n5137, IN2 => n2561, IN3 => RAM_4_43_port, 
                           IN4 => n5126, Q => n1498);
   U1498 : AO22X1 port map( IN1 => RAMDIN1(44), IN2 => n5138, IN3 => 
                           RAM_4_44_port, IN4 => n5125, Q => n1499);
   U1499 : AO22X1 port map( IN1 => n5138, IN2 => RAMDIN1(45), IN3 => 
                           RAM_4_45_port, IN4 => n5125, Q => n1500);
   U1500 : AO22X1 port map( IN1 => RAMDIN1(46), IN2 => n5138, IN3 => 
                           RAM_4_46_port, IN4 => n5125, Q => n1501);
   U1501 : AO22X1 port map( IN1 => n5138, IN2 => RAMDIN1(47), IN3 => 
                           RAM_4_47_port, IN4 => n5125, Q => n1502);
   U1502 : AO22X1 port map( IN1 => n5138, IN2 => n2126, IN3 => RAM_4_48_port, 
                           IN4 => n5125, Q => n1503);
   U1503 : AO22X1 port map( IN1 => n5139, IN2 => RAMDIN1(49), IN3 => 
                           RAM_4_49_port, IN4 => n5125, Q => n1504);
   U1504 : AO22X1 port map( IN1 => n5139, IN2 => RAMDIN1(50), IN3 => 
                           RAM_4_50_port, IN4 => n5125, Q => n1505);
   U1505 : AO22X1 port map( IN1 => n5139, IN2 => RAMDIN1(51), IN3 => 
                           RAM_4_51_port, IN4 => n5125, Q => n1506);
   U1506 : AO22X1 port map( IN1 => n5139, IN2 => n2, IN3 => RAM_4_52_port, IN4 
                           => n5125, Q => n1507);
   U1507 : AO22X1 port map( IN1 => n5139, IN2 => RAMDIN1(53), IN3 => 
                           RAM_4_53_port, IN4 => n5125, Q => n1508);
   U1508 : AO22X1 port map( IN1 => n5140, IN2 => RAMDIN1(54), IN3 => 
                           RAM_4_54_port, IN4 => n5125, Q => n1509);
   U1509 : AO22X1 port map( IN1 => n5140, IN2 => RAMDIN1(55), IN3 => 
                           RAM_4_55_port, IN4 => n5125, Q => n1510);
   U1510 : AO22X1 port map( IN1 => n5140, IN2 => RAMDIN1(56), IN3 => 
                           RAM_4_56_port, IN4 => n5124, Q => n1511);
   U1511 : AO22X1 port map( IN1 => n5140, IN2 => RAMDIN1(57), IN3 => 
                           RAM_4_57_port, IN4 => n5124, Q => n1512);
   U1512 : AO22X1 port map( IN1 => n5140, IN2 => RAMDIN1(58), IN3 => 
                           RAM_4_58_port, IN4 => n5124, Q => n1513);
   U1513 : AO22X1 port map( IN1 => n5141, IN2 => RAMDIN1(59), IN3 => 
                           RAM_4_59_port, IN4 => n5124, Q => n1514);
   U1514 : AO22X1 port map( IN1 => n5141, IN2 => RAMDIN1(60), IN3 => 
                           RAM_4_60_port, IN4 => n5124, Q => n1515);
   U1515 : AO22X1 port map( IN1 => n5141, IN2 => RAMDIN1(61), IN3 => 
                           RAM_4_61_port, IN4 => n5124, Q => n1516);
   U1516 : AO22X1 port map( IN1 => n5141, IN2 => RAMDIN1(62), IN3 => 
                           RAM_4_62_port, IN4 => n5124, Q => n1517);
   U1517 : AO22X1 port map( IN1 => n5141, IN2 => RAMDIN1(63), IN3 => 
                           RAM_4_63_port, IN4 => n5124, Q => n1518);
   U1518 : AO22X1 port map( IN1 => n5142, IN2 => RAMDIN1(64), IN3 => 
                           RAM_4_64_port, IN4 => n5124, Q => n1519);
   U1519 : AO22X1 port map( IN1 => n5142, IN2 => RAMDIN1(65), IN3 => 
                           RAM_4_65_port, IN4 => n5124, Q => n1520);
   U1520 : AO22X1 port map( IN1 => n5142, IN2 => RAMDIN1(66), IN3 => 
                           RAM_4_66_port, IN4 => n5124, Q => n1521);
   U1521 : AO22X1 port map( IN1 => n5142, IN2 => RAMDIN1(67), IN3 => 
                           RAM_4_67_port, IN4 => n5124, Q => n1522);
   U1522 : AO22X1 port map( IN1 => n5142, IN2 => RAMDIN1(68), IN3 => 
                           RAM_4_68_port, IN4 => n5123, Q => n1523);
   U1523 : AO22X1 port map( IN1 => n5143, IN2 => RAMDIN1(69), IN3 => 
                           RAM_4_69_port, IN4 => n5123, Q => n1524);
   U1524 : AO22X1 port map( IN1 => n5143, IN2 => RAMDIN1(70), IN3 => 
                           RAM_4_70_port, IN4 => n5123, Q => n1525);
   U1525 : AO22X1 port map( IN1 => n5143, IN2 => RAMDIN1(71), IN3 => 
                           RAM_4_71_port, IN4 => n5123, Q => n1526);
   U1526 : AO22X1 port map( IN1 => n5143, IN2 => RAMDIN1(72), IN3 => 
                           RAM_4_72_port, IN4 => n5123, Q => n1527);
   U1527 : AO22X1 port map( IN1 => n5143, IN2 => RAMDIN1(73), IN3 => 
                           RAM_4_73_port, IN4 => n5123, Q => n1528);
   U1528 : AO22X1 port map( IN1 => n5144, IN2 => RAMDIN1(74), IN3 => 
                           RAM_4_74_port, IN4 => n5123, Q => n1529);
   U1529 : AO22X1 port map( IN1 => n5144, IN2 => RAMDIN1(75), IN3 => 
                           RAM_4_75_port, IN4 => n5123, Q => n1530);
   U1530 : AO22X1 port map( IN1 => n5144, IN2 => RAMDIN1(76), IN3 => 
                           RAM_4_76_port, IN4 => n5123, Q => n1531);
   U1531 : AO22X1 port map( IN1 => n5144, IN2 => RAMDIN1(77), IN3 => 
                           RAM_4_77_port, IN4 => n5123, Q => n1532);
   U1532 : AO22X1 port map( IN1 => n5144, IN2 => RAMDIN1(78), IN3 => 
                           RAM_4_78_port, IN4 => n5123, Q => n1533);
   U1533 : AO22X1 port map( IN1 => n5145, IN2 => RAMDIN1(79), IN3 => 
                           RAM_4_79_port, IN4 => n5123, Q => n1534);
   U1534 : AO22X1 port map( IN1 => RAMDIN1(80), IN2 => n5145, IN3 => 
                           RAM_4_80_port, IN4 => n5122, Q => n1535);
   U1535 : AO22X1 port map( IN1 => n5145, IN2 => RAMDIN1(81), IN3 => 
                           RAM_4_81_port, IN4 => n5122, Q => n1536);
   U1536 : AO22X1 port map( IN1 => n5145, IN2 => RAMDIN1(82), IN3 => 
                           RAM_4_82_port, IN4 => n5122, Q => n1537);
   U1537 : AO22X1 port map( IN1 => n5145, IN2 => RAMDIN1(83), IN3 => 
                           RAM_4_83_port, IN4 => n5122, Q => n1538);
   U1538 : AO22X1 port map( IN1 => n5146, IN2 => RAMDIN1(84), IN3 => 
                           RAM_4_84_port, IN4 => n5122, Q => n1539);
   U1539 : AO22X1 port map( IN1 => n5146, IN2 => RAMDIN1(85), IN3 => 
                           RAM_4_85_port, IN4 => n5122, Q => n1540);
   U1540 : AO22X1 port map( IN1 => n5146, IN2 => RAMDIN1(86), IN3 => 
                           RAM_4_86_port, IN4 => n5122, Q => n1541);
   U1541 : AO22X1 port map( IN1 => n5146, IN2 => RAMDIN1(87), IN3 => 
                           RAM_4_87_port, IN4 => n5122, Q => n1542);
   U1542 : AO22X1 port map( IN1 => RAMDIN1(88), IN2 => n5146, IN3 => 
                           RAM_4_88_port, IN4 => n5122, Q => n1543);
   U1543 : AO22X1 port map( IN1 => n5147, IN2 => RAMDIN1(89), IN3 => 
                           RAM_4_89_port, IN4 => n5122, Q => n1544);
   U1544 : AO22X1 port map( IN1 => n5147, IN2 => RAMDIN1(90), IN3 => 
                           RAM_4_90_port, IN4 => n5122, Q => n1545);
   U1545 : AO22X1 port map( IN1 => n5147, IN2 => RAMDIN1(91), IN3 => 
                           RAM_4_91_port, IN4 => n5122, Q => n1546);
   U1546 : AO22X1 port map( IN1 => n5147, IN2 => RAMDIN1(92), IN3 => 
                           RAM_4_92_port, IN4 => n5121, Q => n1547);
   U1547 : AO22X1 port map( IN1 => n5147, IN2 => RAMDIN1(93), IN3 => 
                           RAM_4_93_port, IN4 => n5121, Q => n1548);
   U1548 : AO22X1 port map( IN1 => n5148, IN2 => RAMDIN1(94), IN3 => 
                           RAM_4_94_port, IN4 => n5121, Q => n1549);
   U1549 : AO22X1 port map( IN1 => n5148, IN2 => RAMDIN1(95), IN3 => 
                           RAM_4_95_port, IN4 => n5121, Q => n1550);
   U1550 : AO22X1 port map( IN1 => n5148, IN2 => RAMDIN1(96), IN3 => 
                           RAM_4_96_port, IN4 => n5121, Q => n1551);
   U1551 : AO22X1 port map( IN1 => n5148, IN2 => RAMDIN1(97), IN3 => 
                           RAM_4_97_port, IN4 => n5121, Q => n1552);
   U1552 : AO22X1 port map( IN1 => n5148, IN2 => RAMDIN1(98), IN3 => 
                           RAM_4_98_port, IN4 => n5121, Q => n1553);
   U1553 : AO22X1 port map( IN1 => n5149, IN2 => n2503, IN3 => RAM_4_99_port, 
                           IN4 => n5121, Q => n1554);
   U1554 : AO22X1 port map( IN1 => n5149, IN2 => RAMDIN1(100), IN3 => 
                           RAM_4_100_port, IN4 => n5121, Q => n1555);
   U1555 : AO22X1 port map( IN1 => n5149, IN2 => RAMDIN1(101), IN3 => 
                           RAM_4_101_port, IN4 => n5121, Q => n1556);
   U1556 : AO22X1 port map( IN1 => n5149, IN2 => RAMDIN1(102), IN3 => 
                           RAM_4_102_port, IN4 => n5121, Q => n1557);
   U1557 : AO22X1 port map( IN1 => n5149, IN2 => RAMDIN1(103), IN3 => 
                           RAM_4_103_port, IN4 => n5121, Q => n1558);
   U1558 : AO22X1 port map( IN1 => n5150, IN2 => RAMDIN1(104), IN3 => 
                           RAM_4_104_port, IN4 => n5120, Q => n1559);
   U1559 : AO22X1 port map( IN1 => n5150, IN2 => RAMDIN1(105), IN3 => 
                           RAM_4_105_port, IN4 => n5120, Q => n1560);
   U1560 : AO22X1 port map( IN1 => n5150, IN2 => RAMDIN1(106), IN3 => 
                           RAM_4_106_port, IN4 => n5120, Q => n1561);
   U1561 : AO22X1 port map( IN1 => n5150, IN2 => RAMDIN1(107), IN3 => 
                           RAM_4_107_port, IN4 => n5120, Q => n1562);
   U1562 : AO22X1 port map( IN1 => n5150, IN2 => RAMDIN1(108), IN3 => 
                           RAM_4_108_port, IN4 => n5120, Q => n1563);
   U1563 : AO22X1 port map( IN1 => n5151, IN2 => RAMDIN1(109), IN3 => 
                           RAM_4_109_port, IN4 => n5120, Q => n1564);
   U1564 : AO22X1 port map( IN1 => RAMDIN1(110), IN2 => n5151, IN3 => 
                           RAM_4_110_port, IN4 => n5120, Q => n1565);
   U1565 : AO22X1 port map( IN1 => n5151, IN2 => RAMDIN1(111), IN3 => 
                           RAM_4_111_port, IN4 => n5120, Q => n1566);
   U1566 : AO22X1 port map( IN1 => RAMDIN1(112), IN2 => n5151, IN3 => 
                           RAM_4_112_port, IN4 => n5120, Q => n1567);
   U1567 : AO22X1 port map( IN1 => n5151, IN2 => RAMDIN1(113), IN3 => 
                           RAM_4_113_port, IN4 => n5120, Q => n1568);
   U1568 : AO22X1 port map( IN1 => n5152, IN2 => RAMDIN1(114), IN3 => 
                           RAM_4_114_port, IN4 => n5120, Q => n1569);
   U1569 : AO22X1 port map( IN1 => n5152, IN2 => RAMDIN1(115), IN3 => 
                           RAM_4_115_port, IN4 => n5120, Q => n1570);
   U1570 : AO22X1 port map( IN1 => n5152, IN2 => RAMDIN1(116), IN3 => 
                           RAM_4_116_port, IN4 => n5119, Q => n1571);
   U1571 : AO22X1 port map( IN1 => n5152, IN2 => RAMDIN1(117), IN3 => 
                           RAM_4_117_port, IN4 => n5119, Q => n1572);
   U1572 : AO22X1 port map( IN1 => n5152, IN2 => RAMDIN1(118), IN3 => 
                           RAM_4_118_port, IN4 => n5119, Q => n1573);
   U1573 : AO22X1 port map( IN1 => n5153, IN2 => RAMDIN1(119), IN3 => 
                           RAM_4_119_port, IN4 => n5119, Q => n1574);
   U1574 : AO22X1 port map( IN1 => n5153, IN2 => RAMDIN1(120), IN3 => 
                           RAM_4_120_port, IN4 => n5119, Q => n1575);
   U1575 : AO22X1 port map( IN1 => n5153, IN2 => RAMDIN1(121), IN3 => 
                           RAM_4_121_port, IN4 => n5119, Q => n1576);
   U1576 : AO22X1 port map( IN1 => n5153, IN2 => RAMDIN1(122), IN3 => 
                           RAM_4_122_port, IN4 => n5119, Q => n1577);
   U1577 : AO22X1 port map( IN1 => n5153, IN2 => RAMDIN1(123), IN3 => 
                           RAM_4_123_port, IN4 => n5119, Q => n1578);
   U1578 : AO22X1 port map( IN1 => n5154, IN2 => RAMDIN1(124), IN3 => 
                           RAM_4_124_port, IN4 => n5119, Q => n1579);
   U1579 : AO22X1 port map( IN1 => n5154, IN2 => RAMDIN1(125), IN3 => 
                           RAM_4_125_port, IN4 => n5119, Q => n1580);
   U1580 : AO22X1 port map( IN1 => n5154, IN2 => RAMDIN1(126), IN3 => 
                           RAM_4_126_port, IN4 => n5119, Q => n1581);
   U1581 : AO22X1 port map( IN1 => RAMDIN1(127), IN2 => n5154, IN3 => 
                           RAM_4_127_port, IN4 => n5119, Q => n1582);
   U1582 : AO22X1 port map( IN1 => n5092, IN2 => RAMDIN1(0), IN3 => 
                           RAM_3_0_port, IN4 => n5088, Q => n1583);
   U1583 : AO22X1 port map( IN1 => n5091, IN2 => RAMDIN1(1), IN3 => 
                           RAM_3_1_port, IN4 => n5088, Q => n1584);
   U1584 : AO22X1 port map( IN1 => n5089, IN2 => RAMDIN1(2), IN3 => 
                           RAM_3_2_port, IN4 => n5088, Q => n1585);
   U1585 : AO22X1 port map( IN1 => n5089, IN2 => RAMDIN1(3), IN3 => 
                           RAM_3_3_port, IN4 => n5088, Q => n1586);
   U1586 : AO22X1 port map( IN1 => n5111, IN2 => RAMDIN1(4), IN3 => 
                           RAM_3_4_port, IN4 => n5088, Q => n1587);
   U1587 : AO22X1 port map( IN1 => n5112, IN2 => RAMDIN1(5), IN3 => 
                           RAM_3_5_port, IN4 => n5088, Q => n1588);
   U1588 : AO22X1 port map( IN1 => n5111, IN2 => RAMDIN1(6), IN3 => 
                           RAM_3_6_port, IN4 => n5088, Q => n1589);
   U1589 : AO22X1 port map( IN1 => n5112, IN2 => RAMDIN1(7), IN3 => 
                           RAM_3_7_port, IN4 => n5088, Q => n1590);
   U1590 : AO22X1 port map( IN1 => RAMDIN1(8), IN2 => n5110, IN3 => 
                           RAM_3_8_port, IN4 => n5087, Q => n1591);
   U1591 : AO22X1 port map( IN1 => n5112, IN2 => RAMDIN1(9), IN3 => 
                           RAM_3_9_port, IN4 => n5087, Q => n1592);
   U1592 : AO22X1 port map( IN1 => n5111, IN2 => RAMDIN1(10), IN3 => 
                           RAM_3_10_port, IN4 => n5087, Q => n1593);
   U1593 : AO22X1 port map( IN1 => n5110, IN2 => RAMDIN1(11), IN3 => 
                           RAM_3_11_port, IN4 => n5087, Q => n1594);
   U1594 : AO22X1 port map( IN1 => n5112, IN2 => RAMDIN1(12), IN3 => 
                           RAM_3_12_port, IN4 => n5087, Q => n1595);
   U1595 : AO22X1 port map( IN1 => n5110, IN2 => RAMDIN1(13), IN3 => 
                           RAM_3_13_port, IN4 => n5087, Q => n1596);
   U1596 : AO22X1 port map( IN1 => RAMDIN1(14), IN2 => n5091, IN3 => 
                           RAM_3_14_port, IN4 => n5087, Q => n1597);
   U1597 : AO22X1 port map( IN1 => n5091, IN2 => RAMDIN1(15), IN3 => 
                           RAM_3_15_port, IN4 => n5087, Q => n1598);
   U1598 : AO22X1 port map( IN1 => RAMDIN1(16), IN2 => n5091, IN3 => 
                           RAM_3_16_port, IN4 => n5087, Q => n1599);
   U1599 : AO22X1 port map( IN1 => n5091, IN2 => RAMDIN1(17), IN3 => 
                           RAM_3_17_port, IN4 => n5087, Q => n1600);
   U1600 : AO22X1 port map( IN1 => n5091, IN2 => RAMDIN1(18), IN3 => 
                           RAM_3_18_port, IN4 => n5087, Q => n1601);
   U1601 : AO22X1 port map( IN1 => n5092, IN2 => RAMDIN1(19), IN3 => 
                           RAM_3_19_port, IN4 => n5087, Q => n1602);
   U1602 : AO22X1 port map( IN1 => n5092, IN2 => RAMDIN1(20), IN3 => 
                           RAM_3_20_port, IN4 => n5086, Q => n1603);
   U1603 : AO22X1 port map( IN1 => n5092, IN2 => RAMDIN1(21), IN3 => 
                           RAM_3_21_port, IN4 => n5086, Q => n1604);
   U1604 : AO22X1 port map( IN1 => n5092, IN2 => n2103, IN3 => RAM_3_22_port, 
                           IN4 => n5086, Q => n1605);
   U1605 : AO22X1 port map( IN1 => n5092, IN2 => RAMDIN1(23), IN3 => 
                           RAM_3_23_port, IN4 => n5086, Q => n1606);
   U1606 : AO22X1 port map( IN1 => n5093, IN2 => n2200, IN3 => RAM_3_24_port, 
                           IN4 => n5086, Q => n1607);
   U1607 : AO22X1 port map( IN1 => n5093, IN2 => RAMDIN1(25), IN3 => 
                           RAM_3_25_port, IN4 => n5086, Q => n1608);
   U1608 : AO22X1 port map( IN1 => n5093, IN2 => RAMDIN1(26), IN3 => 
                           RAM_3_26_port, IN4 => n5086, Q => n1609);
   U1609 : AO22X1 port map( IN1 => n5093, IN2 => RAMDIN1(27), IN3 => 
                           RAM_3_27_port, IN4 => n5086, Q => n1610);
   U1610 : AO22X1 port map( IN1 => RAMDIN1(28), IN2 => n5093, IN3 => 
                           RAM_3_28_port, IN4 => n5086, Q => n1611);
   U1611 : AO22X1 port map( IN1 => n5094, IN2 => RAMDIN1(29), IN3 => 
                           RAM_3_29_port, IN4 => n5086, Q => n1612);
   U1612 : AO22X1 port map( IN1 => n5094, IN2 => RAMDIN1(30), IN3 => 
                           RAM_3_30_port, IN4 => n5086, Q => n1613);
   U1613 : AO22X1 port map( IN1 => n5094, IN2 => RAMDIN1(31), IN3 => 
                           RAM_3_31_port, IN4 => n5086, Q => n1614);
   U1614 : AO22X1 port map( IN1 => n5094, IN2 => RAMDIN1(32), IN3 => 
                           RAM_3_32_port, IN4 => n5085, Q => n1615);
   U1615 : AO22X1 port map( IN1 => n5094, IN2 => RAMDIN1(33), IN3 => 
                           RAM_3_33_port, IN4 => n5085, Q => n1616);
   U1616 : AO22X1 port map( IN1 => n5092, IN2 => RAMDIN1(34), IN3 => 
                           RAM_3_34_port, IN4 => n5085, Q => n1617);
   U1617 : AO22X1 port map( IN1 => n5094, IN2 => RAMDIN1(35), IN3 => 
                           RAM_3_35_port, IN4 => n5085, Q => n1618);
   U1618 : AO22X1 port map( IN1 => n5093, IN2 => RAMDIN1(36), IN3 => 
                           RAM_3_36_port, IN4 => n5085, Q => n1619);
   U1619 : AO22X1 port map( IN1 => n5094, IN2 => n1, IN3 => RAM_3_37_port, IN4 
                           => n5085, Q => n1620);
   U1620 : AO22X1 port map( IN1 => n5093, IN2 => RAMDIN1(38), IN3 => 
                           RAM_3_38_port, IN4 => n5085, Q => n1621);
   U1621 : AO22X1 port map( IN1 => n5095, IN2 => RAMDIN1(39), IN3 => 
                           RAM_3_39_port, IN4 => n5085, Q => n1622);
   U1622 : AO22X1 port map( IN1 => n5095, IN2 => RAMDIN1(40), IN3 => 
                           RAM_3_40_port, IN4 => n5085, Q => n1623);
   U1623 : AO22X1 port map( IN1 => n5095, IN2 => n2506, IN3 => RAM_3_41_port, 
                           IN4 => n5085, Q => n1624);
   U1624 : AO22X1 port map( IN1 => n5095, IN2 => RAMDIN1(42), IN3 => 
                           RAM_3_42_port, IN4 => n5085, Q => n1625);
   U1625 : AO22X1 port map( IN1 => n5095, IN2 => n2560, IN3 => RAM_3_43_port, 
                           IN4 => n5085, Q => n1626);
   U1626 : AO22X1 port map( IN1 => RAMDIN1(44), IN2 => n5096, IN3 => 
                           RAM_3_44_port, IN4 => n5084, Q => n1627);
   U1627 : AO22X1 port map( IN1 => n5096, IN2 => RAMDIN1(45), IN3 => 
                           RAM_3_45_port, IN4 => n5084, Q => n1628);
   U1628 : AO22X1 port map( IN1 => RAMDIN1(46), IN2 => n5096, IN3 => 
                           RAM_3_46_port, IN4 => n5084, Q => n1629);
   U1629 : AO22X1 port map( IN1 => n5096, IN2 => RAMDIN1(47), IN3 => 
                           RAM_3_47_port, IN4 => n5084, Q => n1630);
   U1630 : AO22X1 port map( IN1 => n5096, IN2 => n2127, IN3 => RAM_3_48_port, 
                           IN4 => n5084, Q => n1631);
   U1631 : AO22X1 port map( IN1 => n5097, IN2 => RAMDIN1(49), IN3 => 
                           RAM_3_49_port, IN4 => n5084, Q => n1632);
   U1632 : AO22X1 port map( IN1 => n5097, IN2 => RAMDIN1(50), IN3 => 
                           RAM_3_50_port, IN4 => n5084, Q => n1633);
   U1633 : AO22X1 port map( IN1 => n5097, IN2 => RAMDIN1(51), IN3 => 
                           RAM_3_51_port, IN4 => n5084, Q => n1634);
   U1634 : AO22X1 port map( IN1 => n5097, IN2 => n2555, IN3 => RAM_3_52_port, 
                           IN4 => n5084, Q => n1635);
   U1635 : AO22X1 port map( IN1 => n5097, IN2 => RAMDIN1(53), IN3 => 
                           RAM_3_53_port, IN4 => n5084, Q => n1636);
   U1636 : AO22X1 port map( IN1 => n5098, IN2 => RAMDIN1(54), IN3 => 
                           RAM_3_54_port, IN4 => n5084, Q => n1637);
   U1637 : AO22X1 port map( IN1 => n5098, IN2 => RAMDIN1(55), IN3 => 
                           RAM_3_55_port, IN4 => n5084, Q => n1638);
   U1638 : AO22X1 port map( IN1 => n5098, IN2 => RAMDIN1(56), IN3 => 
                           RAM_3_56_port, IN4 => n5083, Q => n1639);
   U1639 : AO22X1 port map( IN1 => n5098, IN2 => RAMDIN1(57), IN3 => 
                           RAM_3_57_port, IN4 => n5083, Q => n1640);
   U1640 : AO22X1 port map( IN1 => n5098, IN2 => RAMDIN1(58), IN3 => 
                           RAM_3_58_port, IN4 => n5083, Q => n1641);
   U1641 : AO22X1 port map( IN1 => n5099, IN2 => RAMDIN1(59), IN3 => 
                           RAM_3_59_port, IN4 => n5083, Q => n1642);
   U1642 : AO22X1 port map( IN1 => n5099, IN2 => RAMDIN1(60), IN3 => 
                           RAM_3_60_port, IN4 => n5083, Q => n1643);
   U1643 : AO22X1 port map( IN1 => n5099, IN2 => RAMDIN1(61), IN3 => 
                           RAM_3_61_port, IN4 => n5083, Q => n1644);
   U1644 : AO22X1 port map( IN1 => n5099, IN2 => RAMDIN1(62), IN3 => 
                           RAM_3_62_port, IN4 => n5083, Q => n1645);
   U1645 : AO22X1 port map( IN1 => n5099, IN2 => RAMDIN1(63), IN3 => 
                           RAM_3_63_port, IN4 => n5083, Q => n1646);
   U1646 : AO22X1 port map( IN1 => n5100, IN2 => RAMDIN1(64), IN3 => 
                           RAM_3_64_port, IN4 => n5083, Q => n1647);
   U1647 : AO22X1 port map( IN1 => n5100, IN2 => RAMDIN1(65), IN3 => 
                           RAM_3_65_port, IN4 => n5083, Q => n1648);
   U1648 : AO22X1 port map( IN1 => n5100, IN2 => RAMDIN1(66), IN3 => 
                           RAM_3_66_port, IN4 => n5083, Q => n1649);
   U1649 : AO22X1 port map( IN1 => n5100, IN2 => RAMDIN1(67), IN3 => 
                           RAM_3_67_port, IN4 => n5083, Q => n1650);
   U1650 : AO22X1 port map( IN1 => n5100, IN2 => RAMDIN1(68), IN3 => 
                           RAM_3_68_port, IN4 => n5082, Q => n1651);
   U1651 : AO22X1 port map( IN1 => n5101, IN2 => RAMDIN1(69), IN3 => 
                           RAM_3_69_port, IN4 => n5082, Q => n1652);
   U1652 : AO22X1 port map( IN1 => n5101, IN2 => RAMDIN1(70), IN3 => 
                           RAM_3_70_port, IN4 => n5082, Q => n1653);
   U1653 : AO22X1 port map( IN1 => n5101, IN2 => RAMDIN1(71), IN3 => 
                           RAM_3_71_port, IN4 => n5082, Q => n1654);
   U1654 : AO22X1 port map( IN1 => n5101, IN2 => RAMDIN1(72), IN3 => 
                           RAM_3_72_port, IN4 => n5082, Q => n1655);
   U1655 : AO22X1 port map( IN1 => n5101, IN2 => RAMDIN1(73), IN3 => 
                           RAM_3_73_port, IN4 => n5082, Q => n1656);
   U1656 : AO22X1 port map( IN1 => n5102, IN2 => RAMDIN1(74), IN3 => 
                           RAM_3_74_port, IN4 => n5082, Q => n1657);
   U1657 : AO22X1 port map( IN1 => n5102, IN2 => RAMDIN1(75), IN3 => 
                           RAM_3_75_port, IN4 => n5082, Q => n1658);
   U1658 : AO22X1 port map( IN1 => n5102, IN2 => RAMDIN1(76), IN3 => 
                           RAM_3_76_port, IN4 => n5082, Q => n1659);
   U1659 : AO22X1 port map( IN1 => n5102, IN2 => RAMDIN1(77), IN3 => 
                           RAM_3_77_port, IN4 => n5082, Q => n1660);
   U1660 : AO22X1 port map( IN1 => n5102, IN2 => RAMDIN1(78), IN3 => 
                           RAM_3_78_port, IN4 => n5082, Q => n1661);
   U1661 : AO22X1 port map( IN1 => n5103, IN2 => RAMDIN1(79), IN3 => 
                           RAM_3_79_port, IN4 => n5082, Q => n1662);
   U1662 : AO22X1 port map( IN1 => RAMDIN1(80), IN2 => n5103, IN3 => 
                           RAM_3_80_port, IN4 => n5081, Q => n1663);
   U1663 : AO22X1 port map( IN1 => n5103, IN2 => RAMDIN1(81), IN3 => 
                           RAM_3_81_port, IN4 => n5081, Q => n1664);
   U1664 : AO22X1 port map( IN1 => n5103, IN2 => RAMDIN1(82), IN3 => 
                           RAM_3_82_port, IN4 => n5081, Q => n1665);
   U1665 : AO22X1 port map( IN1 => n5103, IN2 => RAMDIN1(83), IN3 => 
                           RAM_3_83_port, IN4 => n5081, Q => n1666);
   U1666 : AO22X1 port map( IN1 => n5104, IN2 => RAMDIN1(84), IN3 => 
                           RAM_3_84_port, IN4 => n5081, Q => n1667);
   U1667 : AO22X1 port map( IN1 => n5104, IN2 => RAMDIN1(85), IN3 => 
                           RAM_3_85_port, IN4 => n5081, Q => n1668);
   U1668 : AO22X1 port map( IN1 => n5104, IN2 => RAMDIN1(86), IN3 => 
                           RAM_3_86_port, IN4 => n5081, Q => n1669);
   U1669 : AO22X1 port map( IN1 => RAMDIN1(87), IN2 => n5104, IN3 => 
                           RAM_3_87_port, IN4 => n5081, Q => n1670);
   U1670 : AO22X1 port map( IN1 => RAMDIN1(88), IN2 => n5104, IN3 => 
                           RAM_3_88_port, IN4 => n5081, Q => n1671);
   U1671 : AO22X1 port map( IN1 => n5105, IN2 => RAMDIN1(89), IN3 => 
                           RAM_3_89_port, IN4 => n5081, Q => n1672);
   U1672 : AO22X1 port map( IN1 => n5105, IN2 => RAMDIN1(90), IN3 => 
                           RAM_3_90_port, IN4 => n5081, Q => n1673);
   U1673 : AO22X1 port map( IN1 => n5105, IN2 => RAMDIN1(91), IN3 => 
                           RAM_3_91_port, IN4 => n5081, Q => n1674);
   U1674 : AO22X1 port map( IN1 => n5105, IN2 => RAMDIN1(92), IN3 => 
                           RAM_3_92_port, IN4 => n5080, Q => n1675);
   U1675 : AO22X1 port map( IN1 => n5105, IN2 => RAMDIN1(93), IN3 => 
                           RAM_3_93_port, IN4 => n5080, Q => n1676);
   U1676 : AO22X1 port map( IN1 => n5106, IN2 => RAMDIN1(94), IN3 => 
                           RAM_3_94_port, IN4 => n5080, Q => n1677);
   U1677 : AO22X1 port map( IN1 => n5106, IN2 => RAMDIN1(95), IN3 => 
                           RAM_3_95_port, IN4 => n5080, Q => n1678);
   U1678 : AO22X1 port map( IN1 => n5106, IN2 => RAMDIN1(96), IN3 => 
                           RAM_3_96_port, IN4 => n5080, Q => n1679);
   U1679 : AO22X1 port map( IN1 => n5106, IN2 => RAMDIN1(97), IN3 => 
                           RAM_3_97_port, IN4 => n5080, Q => n1680);
   U1680 : AO22X1 port map( IN1 => n5106, IN2 => RAMDIN1(98), IN3 => 
                           RAM_3_98_port, IN4 => n5080, Q => n1681);
   U1681 : AO22X1 port map( IN1 => n5107, IN2 => n2102, IN3 => RAM_3_99_port, 
                           IN4 => n5080, Q => n1682);
   U1682 : AO22X1 port map( IN1 => n5107, IN2 => RAMDIN1(100), IN3 => 
                           RAM_3_100_port, IN4 => n5080, Q => n1683);
   U1683 : AO22X1 port map( IN1 => n5107, IN2 => RAMDIN1(101), IN3 => 
                           RAM_3_101_port, IN4 => n5080, Q => n1684);
   U1684 : AO22X1 port map( IN1 => n5107, IN2 => RAMDIN1(102), IN3 => 
                           RAM_3_102_port, IN4 => n5080, Q => n1685);
   U1685 : AO22X1 port map( IN1 => n5107, IN2 => RAMDIN1(103), IN3 => 
                           RAM_3_103_port, IN4 => n5080, Q => n1686);
   U1686 : AO22X1 port map( IN1 => n5108, IN2 => RAMDIN1(104), IN3 => 
                           RAM_3_104_port, IN4 => n5079, Q => n1687);
   U1687 : AO22X1 port map( IN1 => n5108, IN2 => RAMDIN1(105), IN3 => 
                           RAM_3_105_port, IN4 => n5079, Q => n1688);
   U1688 : AO22X1 port map( IN1 => n5108, IN2 => RAMDIN1(106), IN3 => 
                           RAM_3_106_port, IN4 => n5079, Q => n1689);
   U1689 : AO22X1 port map( IN1 => n5108, IN2 => RAMDIN1(107), IN3 => 
                           RAM_3_107_port, IN4 => n5079, Q => n1690);
   U1690 : AO22X1 port map( IN1 => n5108, IN2 => RAMDIN1(108), IN3 => 
                           RAM_3_108_port, IN4 => n5079, Q => n1691);
   U1691 : AO22X1 port map( IN1 => n5109, IN2 => RAMDIN1(109), IN3 => 
                           RAM_3_109_port, IN4 => n5079, Q => n1692);
   U1692 : AO22X1 port map( IN1 => RAMDIN1(110), IN2 => n5109, IN3 => 
                           RAM_3_110_port, IN4 => n5079, Q => n1693);
   U1693 : AO22X1 port map( IN1 => n5109, IN2 => RAMDIN1(111), IN3 => 
                           RAM_3_111_port, IN4 => n5079, Q => n1694);
   U1694 : AO22X1 port map( IN1 => RAMDIN1(112), IN2 => n5109, IN3 => 
                           RAM_3_112_port, IN4 => n5079, Q => n1695);
   U1695 : AO22X1 port map( IN1 => n5109, IN2 => RAMDIN1(113), IN3 => 
                           RAM_3_113_port, IN4 => n5079, Q => n1696);
   U1696 : AO22X1 port map( IN1 => n5110, IN2 => RAMDIN1(114), IN3 => 
                           RAM_3_114_port, IN4 => n5079, Q => n1697);
   U1697 : AO22X1 port map( IN1 => n5110, IN2 => RAMDIN1(115), IN3 => 
                           RAM_3_115_port, IN4 => n5079, Q => n1698);
   U1698 : AO22X1 port map( IN1 => n5110, IN2 => RAMDIN1(116), IN3 => 
                           RAM_3_116_port, IN4 => n5078, Q => n1699);
   U1699 : AO22X1 port map( IN1 => n5110, IN2 => RAMDIN1(117), IN3 => 
                           RAM_3_117_port, IN4 => n5078, Q => n1700);
   U1700 : AO22X1 port map( IN1 => n5110, IN2 => RAMDIN1(118), IN3 => 
                           RAM_3_118_port, IN4 => n5078, Q => n1701);
   U1701 : AO22X1 port map( IN1 => n5111, IN2 => RAMDIN1(119), IN3 => 
                           RAM_3_119_port, IN4 => n5078, Q => n1702);
   U1702 : AO22X1 port map( IN1 => n5111, IN2 => RAMDIN1(120), IN3 => 
                           RAM_3_120_port, IN4 => n5078, Q => n1703);
   U1703 : AO22X1 port map( IN1 => n5111, IN2 => RAMDIN1(121), IN3 => 
                           RAM_3_121_port, IN4 => n5078, Q => n1704);
   U1704 : AO22X1 port map( IN1 => n5111, IN2 => RAMDIN1(122), IN3 => 
                           RAM_3_122_port, IN4 => n5078, Q => n1705);
   U1705 : AO22X1 port map( IN1 => n5111, IN2 => RAMDIN1(123), IN3 => 
                           RAM_3_123_port, IN4 => n5078, Q => n1706);
   U1706 : AO22X1 port map( IN1 => n5112, IN2 => RAMDIN1(124), IN3 => 
                           RAM_3_124_port, IN4 => n5078, Q => n1707);
   U1707 : AO22X1 port map( IN1 => n5112, IN2 => RAMDIN1(125), IN3 => 
                           RAM_3_125_port, IN4 => n5078, Q => n1708);
   U1708 : AO22X1 port map( IN1 => n5112, IN2 => RAMDIN1(126), IN3 => 
                           RAM_3_126_port, IN4 => n5078, Q => n1709);
   U1709 : AO22X1 port map( IN1 => RAMDIN1(127), IN2 => n5112, IN3 => 
                           RAM_3_127_port, IN4 => n5078, Q => n1710);
   U1710 : AO22X1 port map( IN1 => n5050, IN2 => RAMDIN1(0), IN3 => 
                           RAM_2_0_port, IN4 => n5046, Q => n1711);
   U1711 : AO22X1 port map( IN1 => n5049, IN2 => RAMDIN1(1), IN3 => 
                           RAM_2_1_port, IN4 => n5046, Q => n1712);
   U1712 : AO22X1 port map( IN1 => n5047, IN2 => RAMDIN1(2), IN3 => 
                           RAM_2_2_port, IN4 => n5046, Q => n1713);
   U1713 : AO22X1 port map( IN1 => n5047, IN2 => RAMDIN1(3), IN3 => 
                           RAM_2_3_port, IN4 => n5046, Q => n1714);
   U1714 : AO22X1 port map( IN1 => n5070, IN2 => RAMDIN1(4), IN3 => 
                           RAM_2_4_port, IN4 => n5046, Q => n1715);
   U1715 : AO22X1 port map( IN1 => n5069, IN2 => RAMDIN1(5), IN3 => 
                           RAM_2_5_port, IN4 => n5046, Q => n1716);
   U1716 : AO22X1 port map( IN1 => n5071, IN2 => RAMDIN1(6), IN3 => 
                           RAM_2_6_port, IN4 => n5046, Q => n1717);
   U1717 : AO22X1 port map( IN1 => RAMDIN1(7), IN2 => n5071, IN3 => 
                           RAM_2_7_port, IN4 => n5046, Q => n1718);
   U1718 : AO22X1 port map( IN1 => n5070, IN2 => RAMDIN1(8), IN3 => 
                           RAM_2_8_port, IN4 => n5045, Q => n1719);
   U1719 : AO22X1 port map( IN1 => n5069, IN2 => RAMDIN1(9), IN3 => 
                           RAM_2_9_port, IN4 => n5045, Q => n1720);
   U1720 : AO22X1 port map( IN1 => n5071, IN2 => RAMDIN1(10), IN3 => 
                           RAM_2_10_port, IN4 => n5045, Q => n1721);
   U1721 : AO22X1 port map( IN1 => n5071, IN2 => RAMDIN1(11), IN3 => 
                           RAM_2_11_port, IN4 => n5045, Q => n1722);
   U1722 : AO22X1 port map( IN1 => n5070, IN2 => RAMDIN1(12), IN3 => 
                           RAM_2_12_port, IN4 => n5045, Q => n1723);
   U1723 : AO22X1 port map( IN1 => RAMDIN1(13), IN2 => n5069, IN3 => 
                           RAM_2_13_port, IN4 => n5045, Q => n1724);
   U1724 : AO22X1 port map( IN1 => RAMDIN1(14), IN2 => n5049, IN3 => 
                           RAM_2_14_port, IN4 => n5045, Q => n1725);
   U1725 : AO22X1 port map( IN1 => n5049, IN2 => RAMDIN1(15), IN3 => 
                           RAM_2_15_port, IN4 => n5045, Q => n1726);
   U1726 : AO22X1 port map( IN1 => RAMDIN1(16), IN2 => n5049, IN3 => 
                           RAM_2_16_port, IN4 => n5045, Q => n1727);
   U1727 : AO22X1 port map( IN1 => n5049, IN2 => RAMDIN1(17), IN3 => 
                           RAM_2_17_port, IN4 => n5045, Q => n1728);
   U1728 : AO22X1 port map( IN1 => n5049, IN2 => RAMDIN1(18), IN3 => 
                           RAM_2_18_port, IN4 => n5045, Q => n1729);
   U1729 : AO22X1 port map( IN1 => n5050, IN2 => RAMDIN1(19), IN3 => 
                           RAM_2_19_port, IN4 => n5045, Q => n1730);
   U1730 : AO22X1 port map( IN1 => n5050, IN2 => RAMDIN1(20), IN3 => 
                           RAM_2_20_port, IN4 => n5044, Q => n1731);
   U1731 : AO22X1 port map( IN1 => n5050, IN2 => RAMDIN1(21), IN3 => 
                           RAM_2_21_port, IN4 => n5044, Q => n1732);
   U1732 : AO22X1 port map( IN1 => n5050, IN2 => n2248, IN3 => RAM_2_22_port, 
                           IN4 => n5044, Q => n1733);
   U1733 : AO22X1 port map( IN1 => n5050, IN2 => RAMDIN1(23), IN3 => 
                           RAM_2_23_port, IN4 => n5044, Q => n1734);
   U1734 : AO22X1 port map( IN1 => n5051, IN2 => n2201, IN3 => RAM_2_24_port, 
                           IN4 => n5044, Q => n1735);
   U1735 : AO22X1 port map( IN1 => n5051, IN2 => RAMDIN1(25), IN3 => 
                           RAM_2_25_port, IN4 => n5044, Q => n1736);
   U1736 : AO22X1 port map( IN1 => n5051, IN2 => RAMDIN1(26), IN3 => 
                           RAM_2_26_port, IN4 => n5044, Q => n1737);
   U1737 : AO22X1 port map( IN1 => n5051, IN2 => RAMDIN1(27), IN3 => 
                           RAM_2_27_port, IN4 => n5044, Q => n1738);
   U1738 : AO22X1 port map( IN1 => RAMDIN1(28), IN2 => n5051, IN3 => 
                           RAM_2_28_port, IN4 => n5044, Q => n1739);
   U1739 : AO22X1 port map( IN1 => n5052, IN2 => RAMDIN1(29), IN3 => 
                           RAM_2_29_port, IN4 => n5044, Q => n1740);
   U1740 : AO22X1 port map( IN1 => n5052, IN2 => RAMDIN1(30), IN3 => 
                           RAM_2_30_port, IN4 => n5044, Q => n1741);
   U1741 : AO22X1 port map( IN1 => n5052, IN2 => RAMDIN1(31), IN3 => 
                           RAM_2_31_port, IN4 => n5044, Q => n1742);
   U1742 : AO22X1 port map( IN1 => n5052, IN2 => RAMDIN1(32), IN3 => 
                           RAM_2_32_port, IN4 => n5043, Q => n1743);
   U1743 : AO22X1 port map( IN1 => n5052, IN2 => RAMDIN1(33), IN3 => 
                           RAM_2_33_port, IN4 => n5043, Q => n1744);
   U1744 : AO22X1 port map( IN1 => n5053, IN2 => RAMDIN1(34), IN3 => 
                           RAM_2_34_port, IN4 => n5043, Q => n1745);
   U1745 : AO22X1 port map( IN1 => n5053, IN2 => RAMDIN1(35), IN3 => 
                           RAM_2_35_port, IN4 => n5043, Q => n1746);
   U1746 : AO22X1 port map( IN1 => n5053, IN2 => RAMDIN1(36), IN3 => 
                           RAM_2_36_port, IN4 => n5043, Q => n1747);
   U1747 : AO22X1 port map( IN1 => n5053, IN2 => n1, IN3 => RAM_2_37_port, IN4 
                           => n5043, Q => n1748);
   U1748 : AO22X1 port map( IN1 => n5053, IN2 => RAMDIN1(38), IN3 => 
                           RAM_2_38_port, IN4 => n5043, Q => n1749);
   U1749 : AO22X1 port map( IN1 => n5054, IN2 => RAMDIN1(39), IN3 => 
                           RAM_2_39_port, IN4 => n5043, Q => n1750);
   U1750 : AO22X1 port map( IN1 => n5054, IN2 => RAMDIN1(40), IN3 => 
                           RAM_2_40_port, IN4 => n5043, Q => n1751);
   U1751 : AO22X1 port map( IN1 => n5054, IN2 => n2104, IN3 => RAM_2_41_port, 
                           IN4 => n5043, Q => n1752);
   U1752 : AO22X1 port map( IN1 => n5054, IN2 => RAMDIN1(42), IN3 => 
                           RAM_2_42_port, IN4 => n5043, Q => n1753);
   U1753 : AO22X1 port map( IN1 => n5054, IN2 => n2560, IN3 => RAM_2_43_port, 
                           IN4 => n5043, Q => n1754);
   U1754 : AO22X1 port map( IN1 => RAMDIN1(44), IN2 => n5055, IN3 => 
                           RAM_2_44_port, IN4 => n5042, Q => n1755);
   U1755 : AO22X1 port map( IN1 => n5055, IN2 => RAMDIN1(45), IN3 => 
                           RAM_2_45_port, IN4 => n5042, Q => n1756);
   U1756 : AO22X1 port map( IN1 => RAMDIN1(46), IN2 => n5055, IN3 => 
                           RAM_2_46_port, IN4 => n5042, Q => n1757);
   U1757 : AO22X1 port map( IN1 => n5055, IN2 => RAMDIN1(47), IN3 => 
                           RAM_2_47_port, IN4 => n5042, Q => n1758);
   U1758 : AO22X1 port map( IN1 => n5055, IN2 => n2126, IN3 => RAM_2_48_port, 
                           IN4 => n5042, Q => n1759);
   U1759 : AO22X1 port map( IN1 => n5056, IN2 => RAMDIN1(49), IN3 => 
                           RAM_2_49_port, IN4 => n5042, Q => n1760);
   U1760 : AO22X1 port map( IN1 => n5056, IN2 => RAMDIN1(50), IN3 => 
                           RAM_2_50_port, IN4 => n5042, Q => n1761);
   U1761 : AO22X1 port map( IN1 => n5056, IN2 => RAMDIN1(51), IN3 => 
                           RAM_2_51_port, IN4 => n5042, Q => n1762);
   U1762 : AO22X1 port map( IN1 => n5056, IN2 => n2555, IN3 => RAM_2_52_port, 
                           IN4 => n5042, Q => n1763);
   U1763 : AO22X1 port map( IN1 => n5056, IN2 => RAMDIN1(53), IN3 => 
                           RAM_2_53_port, IN4 => n5042, Q => n1764);
   U1764 : AO22X1 port map( IN1 => n5057, IN2 => RAMDIN1(54), IN3 => 
                           RAM_2_54_port, IN4 => n5042, Q => n1765);
   U1765 : AO22X1 port map( IN1 => n5057, IN2 => RAMDIN1(55), IN3 => 
                           RAM_2_55_port, IN4 => n5042, Q => n1766);
   U1766 : AO22X1 port map( IN1 => n5057, IN2 => RAMDIN1(56), IN3 => 
                           RAM_2_56_port, IN4 => n5041, Q => n1767);
   U1767 : AO22X1 port map( IN1 => n5057, IN2 => RAMDIN1(57), IN3 => 
                           RAM_2_57_port, IN4 => n5041, Q => n1768);
   U1768 : AO22X1 port map( IN1 => n5057, IN2 => RAMDIN1(58), IN3 => 
                           RAM_2_58_port, IN4 => n5041, Q => n1769);
   U1769 : AO22X1 port map( IN1 => n5058, IN2 => RAMDIN1(59), IN3 => 
                           RAM_2_59_port, IN4 => n5041, Q => n1770);
   U1770 : AO22X1 port map( IN1 => n5058, IN2 => RAMDIN1(60), IN3 => 
                           RAM_2_60_port, IN4 => n5041, Q => n1771);
   U1771 : AO22X1 port map( IN1 => n5058, IN2 => RAMDIN1(61), IN3 => 
                           RAM_2_61_port, IN4 => n5041, Q => n1772);
   U1772 : AO22X1 port map( IN1 => n5058, IN2 => RAMDIN1(62), IN3 => 
                           RAM_2_62_port, IN4 => n5041, Q => n1773);
   U1773 : AO22X1 port map( IN1 => n5058, IN2 => RAMDIN1(63), IN3 => 
                           RAM_2_63_port, IN4 => n5041, Q => n1774);
   U1774 : AO22X1 port map( IN1 => n5059, IN2 => RAMDIN1(64), IN3 => 
                           RAM_2_64_port, IN4 => n5041, Q => n1775);
   U1775 : AO22X1 port map( IN1 => n5059, IN2 => RAMDIN1(65), IN3 => 
                           RAM_2_65_port, IN4 => n5041, Q => n1776);
   U1776 : AO22X1 port map( IN1 => n5059, IN2 => RAMDIN1(66), IN3 => 
                           RAM_2_66_port, IN4 => n5041, Q => n1777);
   U1777 : AO22X1 port map( IN1 => n5059, IN2 => RAMDIN1(67), IN3 => 
                           RAM_2_67_port, IN4 => n5041, Q => n1778);
   U1778 : AO22X1 port map( IN1 => n5059, IN2 => RAMDIN1(68), IN3 => 
                           RAM_2_68_port, IN4 => n5040, Q => n1779);
   U1779 : AO22X1 port map( IN1 => n5060, IN2 => RAMDIN1(69), IN3 => 
                           RAM_2_69_port, IN4 => n5040, Q => n1780);
   U1780 : AO22X1 port map( IN1 => n5060, IN2 => RAMDIN1(70), IN3 => 
                           RAM_2_70_port, IN4 => n5040, Q => n1781);
   U1781 : AO22X1 port map( IN1 => n5060, IN2 => RAMDIN1(71), IN3 => 
                           RAM_2_71_port, IN4 => n5040, Q => n1782);
   U1782 : AO22X1 port map( IN1 => n5060, IN2 => RAMDIN1(72), IN3 => 
                           RAM_2_72_port, IN4 => n5040, Q => n1783);
   U1783 : AO22X1 port map( IN1 => n5060, IN2 => RAMDIN1(73), IN3 => 
                           RAM_2_73_port, IN4 => n5040, Q => n1784);
   U1784 : AO22X1 port map( IN1 => n5061, IN2 => RAMDIN1(74), IN3 => 
                           RAM_2_74_port, IN4 => n5040, Q => n1785);
   U1785 : AO22X1 port map( IN1 => n5061, IN2 => RAMDIN1(75), IN3 => 
                           RAM_2_75_port, IN4 => n5040, Q => n1786);
   U1786 : AO22X1 port map( IN1 => RAMDIN1(76), IN2 => n5061, IN3 => 
                           RAM_2_76_port, IN4 => n5040, Q => n1787);
   U1787 : AO22X1 port map( IN1 => n5061, IN2 => RAMDIN1(77), IN3 => 
                           RAM_2_77_port, IN4 => n5040, Q => n1788);
   U1788 : AO22X1 port map( IN1 => n5061, IN2 => RAMDIN1(78), IN3 => 
                           RAM_2_78_port, IN4 => n5040, Q => n1789);
   U1789 : AO22X1 port map( IN1 => RAMDIN1(79), IN2 => n5062, IN3 => 
                           RAM_2_79_port, IN4 => n5040, Q => n1790);
   U1790 : AO22X1 port map( IN1 => RAMDIN1(80), IN2 => n5062, IN3 => 
                           RAM_2_80_port, IN4 => n5039, Q => n1791);
   U1791 : AO22X1 port map( IN1 => n5062, IN2 => RAMDIN1(81), IN3 => 
                           RAM_2_81_port, IN4 => n5039, Q => n1792);
   U1792 : AO22X1 port map( IN1 => n5062, IN2 => RAMDIN1(82), IN3 => 
                           RAM_2_82_port, IN4 => n5039, Q => n1793);
   U1793 : AO22X1 port map( IN1 => n5062, IN2 => RAMDIN1(83), IN3 => 
                           RAM_2_83_port, IN4 => n5039, Q => n1794);
   U1794 : AO22X1 port map( IN1 => n5063, IN2 => RAMDIN1(84), IN3 => 
                           RAM_2_84_port, IN4 => n5039, Q => n1795);
   U1795 : AO22X1 port map( IN1 => n5063, IN2 => RAMDIN1(85), IN3 => 
                           RAM_2_85_port, IN4 => n5039, Q => n1796);
   U1796 : AO22X1 port map( IN1 => n5063, IN2 => RAMDIN1(86), IN3 => 
                           RAM_2_86_port, IN4 => n5039, Q => n1797);
   U1797 : AO22X1 port map( IN1 => RAMDIN1(87), IN2 => n5063, IN3 => 
                           RAM_2_87_port, IN4 => n5039, Q => n1798);
   U1798 : AO22X1 port map( IN1 => RAMDIN1(88), IN2 => n5063, IN3 => 
                           RAM_2_88_port, IN4 => n5039, Q => n1799);
   U1799 : AO22X1 port map( IN1 => n5064, IN2 => RAMDIN1(89), IN3 => 
                           RAM_2_89_port, IN4 => n5039, Q => n1800);
   U1800 : AO22X1 port map( IN1 => n5064, IN2 => RAMDIN1(90), IN3 => 
                           RAM_2_90_port, IN4 => n5039, Q => n1801);
   U1801 : AO22X1 port map( IN1 => n5064, IN2 => RAMDIN1(91), IN3 => 
                           RAM_2_91_port, IN4 => n5039, Q => n1802);
   U1802 : AO22X1 port map( IN1 => n5064, IN2 => RAMDIN1(92), IN3 => 
                           RAM_2_92_port, IN4 => n5038, Q => n1803);
   U1803 : AO22X1 port map( IN1 => n5064, IN2 => RAMDIN1(93), IN3 => 
                           RAM_2_93_port, IN4 => n5038, Q => n1804);
   U1804 : AO22X1 port map( IN1 => n5065, IN2 => RAMDIN1(94), IN3 => 
                           RAM_2_94_port, IN4 => n5038, Q => n1805);
   U1805 : AO22X1 port map( IN1 => n5065, IN2 => RAMDIN1(95), IN3 => 
                           RAM_2_95_port, IN4 => n5038, Q => n1806);
   U1806 : AO22X1 port map( IN1 => n5065, IN2 => RAMDIN1(96), IN3 => 
                           RAM_2_96_port, IN4 => n5038, Q => n1807);
   U1807 : AO22X1 port map( IN1 => n5065, IN2 => RAMDIN1(97), IN3 => 
                           RAM_2_97_port, IN4 => n5038, Q => n1808);
   U1808 : AO22X1 port map( IN1 => n5065, IN2 => RAMDIN1(98), IN3 => 
                           RAM_2_98_port, IN4 => n5038, Q => n1809);
   U1809 : AO22X1 port map( IN1 => n5066, IN2 => n2502, IN3 => RAM_2_99_port, 
                           IN4 => n5038, Q => n1810);
   U1810 : AO22X1 port map( IN1 => n5066, IN2 => RAMDIN1(100), IN3 => 
                           RAM_2_100_port, IN4 => n5038, Q => n1811);
   U1811 : AO22X1 port map( IN1 => n5066, IN2 => RAMDIN1(101), IN3 => 
                           RAM_2_101_port, IN4 => n5038, Q => n1812);
   U1812 : AO22X1 port map( IN1 => n5066, IN2 => RAMDIN1(102), IN3 => 
                           RAM_2_102_port, IN4 => n5038, Q => n1813);
   U1813 : AO22X1 port map( IN1 => n5066, IN2 => RAMDIN1(103), IN3 => 
                           RAM_2_103_port, IN4 => n5038, Q => n1814);
   U1814 : AO22X1 port map( IN1 => n5067, IN2 => RAMDIN1(104), IN3 => 
                           RAM_2_104_port, IN4 => n5037, Q => n1815);
   U1815 : AO22X1 port map( IN1 => n5067, IN2 => RAMDIN1(105), IN3 => 
                           RAM_2_105_port, IN4 => n5037, Q => n1816);
   U1816 : AO22X1 port map( IN1 => n5067, IN2 => RAMDIN1(106), IN3 => 
                           RAM_2_106_port, IN4 => n5037, Q => n1817);
   U1817 : AO22X1 port map( IN1 => n5067, IN2 => RAMDIN1(107), IN3 => 
                           RAM_2_107_port, IN4 => n5037, Q => n1818);
   U1818 : AO22X1 port map( IN1 => n5067, IN2 => RAMDIN1(108), IN3 => 
                           RAM_2_108_port, IN4 => n5037, Q => n1819);
   U1819 : AO22X1 port map( IN1 => n5068, IN2 => RAMDIN1(109), IN3 => 
                           RAM_2_109_port, IN4 => n5037, Q => n1820);
   U1820 : AO22X1 port map( IN1 => RAMDIN1(110), IN2 => n5068, IN3 => 
                           RAM_2_110_port, IN4 => n5037, Q => n1821);
   U1821 : AO22X1 port map( IN1 => n5068, IN2 => RAMDIN1(111), IN3 => 
                           RAM_2_111_port, IN4 => n5037, Q => n1822);
   U1822 : AO22X1 port map( IN1 => RAMDIN1(112), IN2 => n5068, IN3 => 
                           RAM_2_112_port, IN4 => n5037, Q => n1823);
   U1823 : AO22X1 port map( IN1 => n5068, IN2 => RAMDIN1(113), IN3 => 
                           RAM_2_113_port, IN4 => n5037, Q => n1824);
   U1824 : AO22X1 port map( IN1 => n5069, IN2 => RAMDIN1(114), IN3 => 
                           RAM_2_114_port, IN4 => n5037, Q => n1825);
   U1825 : AO22X1 port map( IN1 => n5069, IN2 => RAMDIN1(115), IN3 => 
                           RAM_2_115_port, IN4 => n5037, Q => n1826);
   U1826 : AO22X1 port map( IN1 => n5069, IN2 => RAMDIN1(116), IN3 => 
                           RAM_2_116_port, IN4 => n5036, Q => n1827);
   U1827 : AO22X1 port map( IN1 => n5069, IN2 => RAMDIN1(117), IN3 => 
                           RAM_2_117_port, IN4 => n5036, Q => n1828);
   U1828 : AO22X1 port map( IN1 => n5069, IN2 => RAMDIN1(118), IN3 => 
                           RAM_2_118_port, IN4 => n5036, Q => n1829);
   U1829 : AO22X1 port map( IN1 => n5070, IN2 => RAMDIN1(119), IN3 => 
                           RAM_2_119_port, IN4 => n5036, Q => n1830);
   U1830 : AO22X1 port map( IN1 => RAMDIN1(120), IN2 => n5070, IN3 => 
                           RAM_2_120_port, IN4 => n5036, Q => n1831);
   U1831 : AO22X1 port map( IN1 => n5070, IN2 => RAMDIN1(121), IN3 => 
                           RAM_2_121_port, IN4 => n5036, Q => n1832);
   U1832 : AO22X1 port map( IN1 => n5070, IN2 => RAMDIN1(122), IN3 => 
                           RAM_2_122_port, IN4 => n5036, Q => n1833);
   U1833 : AO22X1 port map( IN1 => n5070, IN2 => RAMDIN1(123), IN3 => 
                           RAM_2_123_port, IN4 => n5036, Q => n1834);
   U1834 : AO22X1 port map( IN1 => n5071, IN2 => RAMDIN1(124), IN3 => 
                           RAM_2_124_port, IN4 => n5036, Q => n1835);
   U1835 : AO22X1 port map( IN1 => n5071, IN2 => RAMDIN1(125), IN3 => 
                           RAM_2_125_port, IN4 => n5036, Q => n1836);
   U1836 : AO22X1 port map( IN1 => n5071, IN2 => RAMDIN1(126), IN3 => 
                           RAM_2_126_port, IN4 => n5036, Q => n1837);
   U1837 : AO22X1 port map( IN1 => RAMDIN1(127), IN2 => n5071, IN3 => 
                           RAM_2_127_port, IN4 => n5036, Q => n1838);
   U1838 : AO22X1 port map( IN1 => n5010, IN2 => RAMDIN1(0), IN3 => 
                           RAM_1_0_port, IN4 => n5004, Q => n1839);
   U1839 : AO22X1 port map( IN1 => n5009, IN2 => RAMDIN1(1), IN3 => 
                           RAM_1_1_port, IN4 => n5004, Q => n1840);
   U1840 : AO22X1 port map( IN1 => n5006, IN2 => RAMDIN1(2), IN3 => 
                           RAM_1_2_port, IN4 => n5004, Q => n1841);
   U1841 : AO22X1 port map( IN1 => n5006, IN2 => RAMDIN1(3), IN3 => 
                           RAM_1_3_port, IN4 => n5004, Q => n1842);
   U1842 : AO22X1 port map( IN1 => n5028, IN2 => RAMDIN1(4), IN3 => 
                           RAM_1_4_port, IN4 => n5004, Q => n1843);
   U1843 : AO22X1 port map( IN1 => n5027, IN2 => RAMDIN1(5), IN3 => 
                           RAM_1_5_port, IN4 => n5004, Q => n1844);
   U1844 : AO22X1 port map( IN1 => n5029, IN2 => RAMDIN1(6), IN3 => 
                           RAM_1_6_port, IN4 => n5004, Q => n1845);
   U1845 : AO22X1 port map( IN1 => n5028, IN2 => RAMDIN1(7), IN3 => 
                           RAM_1_7_port, IN4 => n5004, Q => n1846);
   U1846 : AO22X1 port map( IN1 => RAMDIN1(8), IN2 => n5029, IN3 => 
                           RAM_1_8_port, IN4 => n5003, Q => n1847);
   U1847 : AO22X1 port map( IN1 => n5027, IN2 => RAMDIN1(9), IN3 => 
                           RAM_1_9_port, IN4 => n5003, Q => n1848);
   U1848 : AO22X1 port map( IN1 => n5028, IN2 => RAMDIN1(10), IN3 => 
                           RAM_1_10_port, IN4 => n5003, Q => n1849);
   U1849 : AO22X1 port map( IN1 => n5027, IN2 => RAMDIN1(11), IN3 => 
                           RAM_1_11_port, IN4 => n5003, Q => n1850);
   U1850 : AO22X1 port map( IN1 => n5029, IN2 => RAMDIN1(12), IN3 => 
                           RAM_1_12_port, IN4 => n5003, Q => n1851);
   U1851 : AO22X1 port map( IN1 => n5029, IN2 => RAMDIN1(13), IN3 => 
                           RAM_1_13_port, IN4 => n5003, Q => n1852);
   U1852 : AO22X1 port map( IN1 => RAMDIN1(14), IN2 => n5007, IN3 => 
                           RAM_1_14_port, IN4 => n5003, Q => n1853);
   U1853 : AO22X1 port map( IN1 => n5007, IN2 => RAMDIN1(15), IN3 => 
                           RAM_1_15_port, IN4 => n5003, Q => n1854);
   U1854 : AO22X1 port map( IN1 => RAMDIN1(16), IN2 => n5007, IN3 => 
                           RAM_1_16_port, IN4 => n5003, Q => n1855);
   U1855 : AO22X1 port map( IN1 => n5007, IN2 => RAMDIN1(17), IN3 => 
                           RAM_1_17_port, IN4 => n5003, Q => n1856);
   U1856 : AO22X1 port map( IN1 => n5007, IN2 => RAMDIN1(18), IN3 => 
                           RAM_1_18_port, IN4 => n5003, Q => n1857);
   U1857 : AO22X1 port map( IN1 => n5008, IN2 => RAMDIN1(19), IN3 => 
                           RAM_1_19_port, IN4 => n5003, Q => n1858);
   U1858 : AO22X1 port map( IN1 => n5008, IN2 => RAMDIN1(20), IN3 => 
                           RAM_1_20_port, IN4 => n5002, Q => n1859);
   U1859 : AO22X1 port map( IN1 => n5008, IN2 => RAMDIN1(21), IN3 => 
                           RAM_1_21_port, IN4 => n5002, Q => n1860);
   U1860 : AO22X1 port map( IN1 => n5008, IN2 => n2249, IN3 => RAM_1_22_port, 
                           IN4 => n5002, Q => n1861);
   U1861 : AO22X1 port map( IN1 => RAMDIN1(23), IN2 => n5008, IN3 => 
                           RAM_1_23_port, IN4 => n5002, Q => n1862);
   U1862 : AO22X1 port map( IN1 => n5009, IN2 => n2200, IN3 => RAM_1_24_port, 
                           IN4 => n5002, Q => n1863);
   U1863 : AO22X1 port map( IN1 => n5009, IN2 => RAMDIN1(25), IN3 => 
                           RAM_1_25_port, IN4 => n5002, Q => n1864);
   U1864 : AO22X1 port map( IN1 => n5009, IN2 => RAMDIN1(26), IN3 => 
                           RAM_1_26_port, IN4 => n5002, Q => n1865);
   U1865 : AO22X1 port map( IN1 => n5009, IN2 => RAMDIN1(27), IN3 => 
                           RAM_1_27_port, IN4 => n5002, Q => n1866);
   U1866 : AO22X1 port map( IN1 => RAMDIN1(28), IN2 => n5009, IN3 => 
                           RAM_1_28_port, IN4 => n5002, Q => n1867);
   U1867 : AO22X1 port map( IN1 => n5010, IN2 => RAMDIN1(29), IN3 => 
                           RAM_1_29_port, IN4 => n5002, Q => n1868);
   U1868 : AO22X1 port map( IN1 => n5010, IN2 => RAMDIN1(30), IN3 => 
                           RAM_1_30_port, IN4 => n5002, Q => n1869);
   U1869 : AO22X1 port map( IN1 => n5010, IN2 => RAMDIN1(31), IN3 => 
                           RAM_1_31_port, IN4 => n5002, Q => n1870);
   U1870 : AO22X1 port map( IN1 => n5010, IN2 => RAMDIN1(32), IN3 => 
                           RAM_1_32_port, IN4 => n5001, Q => n1871);
   U1871 : AO22X1 port map( IN1 => n5010, IN2 => RAMDIN1(33), IN3 => 
                           RAM_1_33_port, IN4 => n5001, Q => n1872);
   U1872 : AO22X1 port map( IN1 => n5011, IN2 => RAMDIN1(34), IN3 => 
                           RAM_1_34_port, IN4 => n5001, Q => n1873);
   U1873 : AO22X1 port map( IN1 => n5011, IN2 => RAMDIN1(35), IN3 => 
                           RAM_1_35_port, IN4 => n5001, Q => n1874);
   U1874 : AO22X1 port map( IN1 => n5011, IN2 => RAMDIN1(36), IN3 => 
                           RAM_1_36_port, IN4 => n5001, Q => n1875);
   U1875 : AO22X1 port map( IN1 => n5011, IN2 => n2559, IN3 => RAM_1_37_port, 
                           IN4 => n5001, Q => n1876);
   U1876 : AO22X1 port map( IN1 => n5011, IN2 => RAMDIN1(38), IN3 => 
                           RAM_1_38_port, IN4 => n5001, Q => n1877);
   U1877 : AO22X1 port map( IN1 => n5012, IN2 => RAMDIN1(39), IN3 => 
                           RAM_1_39_port, IN4 => n5001, Q => n1878);
   U1878 : AO22X1 port map( IN1 => RAMDIN1(40), IN2 => n5012, IN3 => 
                           RAM_1_40_port, IN4 => n5001, Q => n1879);
   U1879 : AO22X1 port map( IN1 => n5012, IN2 => n2506, IN3 => RAM_1_41_port, 
                           IN4 => n5001, Q => n1880);
   U1880 : AO22X1 port map( IN1 => n5012, IN2 => RAMDIN1(42), IN3 => 
                           RAM_1_42_port, IN4 => n5001, Q => n1881);
   U1881 : AO22X1 port map( IN1 => n5012, IN2 => n2561, IN3 => RAM_1_43_port, 
                           IN4 => n5001, Q => n1882);
   U1882 : AO22X1 port map( IN1 => n5013, IN2 => RAMDIN1(44), IN3 => 
                           RAM_1_44_port, IN4 => n5000, Q => n1883);
   U1883 : AO22X1 port map( IN1 => n5013, IN2 => RAMDIN1(45), IN3 => 
                           RAM_1_45_port, IN4 => n5000, Q => n1884);
   U1884 : AO22X1 port map( IN1 => RAMDIN1(46), IN2 => n5013, IN3 => 
                           RAM_1_46_port, IN4 => n5000, Q => n1885);
   U1885 : AO22X1 port map( IN1 => n5013, IN2 => RAMDIN1(47), IN3 => 
                           RAM_1_47_port, IN4 => n5000, Q => n1886);
   U1886 : AO22X1 port map( IN1 => n5013, IN2 => n2557, IN3 => RAM_1_48_port, 
                           IN4 => n5000, Q => n1887);
   U1887 : AO22X1 port map( IN1 => n5014, IN2 => RAMDIN1(49), IN3 => 
                           RAM_1_49_port, IN4 => n5000, Q => n1888);
   U1888 : AO22X1 port map( IN1 => n5014, IN2 => RAMDIN1(50), IN3 => 
                           RAM_1_50_port, IN4 => n5000, Q => n1889);
   U1889 : AO22X1 port map( IN1 => n5014, IN2 => RAMDIN1(51), IN3 => 
                           RAM_1_51_port, IN4 => n5000, Q => n1890);
   U1890 : AO22X1 port map( IN1 => n5014, IN2 => n2556, IN3 => RAM_1_52_port, 
                           IN4 => n5000, Q => n1891);
   U1891 : AO22X1 port map( IN1 => n5014, IN2 => RAMDIN1(53), IN3 => 
                           RAM_1_53_port, IN4 => n5000, Q => n1892);
   U1892 : AO22X1 port map( IN1 => n5015, IN2 => RAMDIN1(54), IN3 => 
                           RAM_1_54_port, IN4 => n5000, Q => n1893);
   U1893 : AO22X1 port map( IN1 => n5015, IN2 => RAMDIN1(55), IN3 => 
                           RAM_1_55_port, IN4 => n5000, Q => n1894);
   U1894 : AO22X1 port map( IN1 => n5015, IN2 => RAMDIN1(56), IN3 => 
                           RAM_1_56_port, IN4 => n4999, Q => n1895);
   U1895 : AO22X1 port map( IN1 => n5015, IN2 => RAMDIN1(57), IN3 => 
                           RAM_1_57_port, IN4 => n4999, Q => n1896);
   U1896 : AO22X1 port map( IN1 => n5015, IN2 => RAMDIN1(58), IN3 => 
                           RAM_1_58_port, IN4 => n4999, Q => n1897);
   U1897 : AO22X1 port map( IN1 => n5016, IN2 => RAMDIN1(59), IN3 => 
                           RAM_1_59_port, IN4 => n4999, Q => n1898);
   U1898 : AO22X1 port map( IN1 => n5016, IN2 => RAMDIN1(60), IN3 => 
                           RAM_1_60_port, IN4 => n4999, Q => n1899);
   U1899 : AO22X1 port map( IN1 => n5016, IN2 => RAMDIN1(61), IN3 => 
                           RAM_1_61_port, IN4 => n4999, Q => n1900);
   U1900 : AO22X1 port map( IN1 => n5016, IN2 => RAMDIN1(62), IN3 => 
                           RAM_1_62_port, IN4 => n4999, Q => n1901);
   U1901 : AO22X1 port map( IN1 => n5016, IN2 => RAMDIN1(63), IN3 => 
                           RAM_1_63_port, IN4 => n4999, Q => n1902);
   U1902 : AO22X1 port map( IN1 => n5017, IN2 => RAMDIN1(64), IN3 => 
                           RAM_1_64_port, IN4 => n4999, Q => n1903);
   U1903 : AO22X1 port map( IN1 => n5017, IN2 => RAMDIN1(65), IN3 => 
                           RAM_1_65_port, IN4 => n4999, Q => n1904);
   U1904 : AO22X1 port map( IN1 => n5017, IN2 => RAMDIN1(66), IN3 => 
                           RAM_1_66_port, IN4 => n4999, Q => n1905);
   U1905 : AO22X1 port map( IN1 => n5017, IN2 => RAMDIN1(67), IN3 => 
                           RAM_1_67_port, IN4 => n4999, Q => n1906);
   U1906 : AO22X1 port map( IN1 => RAMDIN1(68), IN2 => n5017, IN3 => 
                           RAM_1_68_port, IN4 => n4998, Q => n1907);
   U1907 : AO22X1 port map( IN1 => n5018, IN2 => RAMDIN1(69), IN3 => 
                           RAM_1_69_port, IN4 => n4998, Q => n1908);
   U1908 : AO22X1 port map( IN1 => n5018, IN2 => RAMDIN1(70), IN3 => 
                           RAM_1_70_port, IN4 => n4998, Q => n1909);
   U1909 : AO22X1 port map( IN1 => n5018, IN2 => RAMDIN1(71), IN3 => 
                           RAM_1_71_port, IN4 => n4998, Q => n1910);
   U1910 : AO22X1 port map( IN1 => n5018, IN2 => RAMDIN1(72), IN3 => 
                           RAM_1_72_port, IN4 => n4998, Q => n1911);
   U1911 : AO22X1 port map( IN1 => RAMDIN1(73), IN2 => n5018, IN3 => 
                           RAM_1_73_port, IN4 => n4998, Q => n1912);
   U1912 : AO22X1 port map( IN1 => n5019, IN2 => RAMDIN1(74), IN3 => 
                           RAM_1_74_port, IN4 => n4998, Q => n1913);
   U1913 : AO22X1 port map( IN1 => n5019, IN2 => RAMDIN1(75), IN3 => 
                           RAM_1_75_port, IN4 => n4998, Q => n1914);
   U1914 : AO22X1 port map( IN1 => n5019, IN2 => RAMDIN1(76), IN3 => 
                           RAM_1_76_port, IN4 => n4998, Q => n1915);
   U1915 : AO22X1 port map( IN1 => n5019, IN2 => RAMDIN1(77), IN3 => 
                           RAM_1_77_port, IN4 => n4998, Q => n1916);
   U1916 : AO22X1 port map( IN1 => RAMDIN1(78), IN2 => n5019, IN3 => 
                           RAM_1_78_port, IN4 => n4998, Q => n1917);
   U1917 : AO22X1 port map( IN1 => n5020, IN2 => RAMDIN1(79), IN3 => 
                           RAM_1_79_port, IN4 => n4998, Q => n1918);
   U1918 : AO22X1 port map( IN1 => RAMDIN1(80), IN2 => n5020, IN3 => 
                           RAM_1_80_port, IN4 => n4997, Q => n1919);
   U1919 : AO22X1 port map( IN1 => n5020, IN2 => RAMDIN1(81), IN3 => 
                           RAM_1_81_port, IN4 => n4997, Q => n1920);
   U1920 : AO22X1 port map( IN1 => n5020, IN2 => RAMDIN1(82), IN3 => 
                           RAM_1_82_port, IN4 => n4997, Q => n1921);
   U1921 : AO22X1 port map( IN1 => RAMDIN1(83), IN2 => n5020, IN3 => 
                           RAM_1_83_port, IN4 => n4997, Q => n1922);
   U1922 : AO22X1 port map( IN1 => n5021, IN2 => RAMDIN1(84), IN3 => 
                           RAM_1_84_port, IN4 => n4997, Q => n1923);
   U1923 : AO22X1 port map( IN1 => RAMDIN1(85), IN2 => n5021, IN3 => 
                           RAM_1_85_port, IN4 => n4997, Q => n1924);
   U1924 : AO22X1 port map( IN1 => n5021, IN2 => RAMDIN1(86), IN3 => 
                           RAM_1_86_port, IN4 => n4997, Q => n1925);
   U1925 : AO22X1 port map( IN1 => n5021, IN2 => RAMDIN1(87), IN3 => 
                           RAM_1_87_port, IN4 => n4997, Q => n1926);
   U1926 : AO22X1 port map( IN1 => RAMDIN1(88), IN2 => n5021, IN3 => 
                           RAM_1_88_port, IN4 => n4997, Q => n1927);
   U1927 : AO22X1 port map( IN1 => n5022, IN2 => RAMDIN1(89), IN3 => 
                           RAM_1_89_port, IN4 => n4997, Q => n1928);
   U1928 : AO22X1 port map( IN1 => n5022, IN2 => RAMDIN1(90), IN3 => 
                           RAM_1_90_port, IN4 => n4997, Q => n1929);
   U1929 : AO22X1 port map( IN1 => n5022, IN2 => RAMDIN1(91), IN3 => 
                           RAM_1_91_port, IN4 => n4997, Q => n1930);
   U1930 : AO22X1 port map( IN1 => n5022, IN2 => RAMDIN1(92), IN3 => 
                           RAM_1_92_port, IN4 => n4996, Q => n1931);
   U1931 : AO22X1 port map( IN1 => n5022, IN2 => RAMDIN1(93), IN3 => 
                           RAM_1_93_port, IN4 => n4996, Q => n1932);
   U1932 : AO22X1 port map( IN1 => n5023, IN2 => RAMDIN1(94), IN3 => 
                           RAM_1_94_port, IN4 => n4996, Q => n1933);
   U1933 : AO22X1 port map( IN1 => n5023, IN2 => RAMDIN1(95), IN3 => 
                           RAM_1_95_port, IN4 => n4996, Q => n1934);
   U1934 : AO22X1 port map( IN1 => n5023, IN2 => RAMDIN1(96), IN3 => 
                           RAM_1_96_port, IN4 => n4996, Q => n1935);
   U1935 : AO22X1 port map( IN1 => n5023, IN2 => RAMDIN1(97), IN3 => 
                           RAM_1_97_port, IN4 => n4996, Q => n1936);
   U1936 : AO22X1 port map( IN1 => n5023, IN2 => RAMDIN1(98), IN3 => 
                           RAM_1_98_port, IN4 => n4996, Q => n1937);
   U1937 : AO22X1 port map( IN1 => n5024, IN2 => n2503, IN3 => RAM_1_99_port, 
                           IN4 => n4996, Q => n1938);
   U1938 : AO22X1 port map( IN1 => n5024, IN2 => RAMDIN1(100), IN3 => 
                           RAM_1_100_port, IN4 => n4996, Q => n1939);
   U1939 : AO22X1 port map( IN1 => n5024, IN2 => RAMDIN1(101), IN3 => 
                           RAM_1_101_port, IN4 => n4996, Q => n1940);
   U1940 : AO22X1 port map( IN1 => n5024, IN2 => RAMDIN1(102), IN3 => 
                           RAM_1_102_port, IN4 => n4996, Q => n1941);
   U1941 : AO22X1 port map( IN1 => n5024, IN2 => RAMDIN1(103), IN3 => 
                           RAM_1_103_port, IN4 => n4996, Q => n1942);
   U1942 : AO22X1 port map( IN1 => n5025, IN2 => RAMDIN1(104), IN3 => 
                           RAM_1_104_port, IN4 => n4995, Q => n1943);
   U1943 : AO22X1 port map( IN1 => n5025, IN2 => RAMDIN1(105), IN3 => 
                           RAM_1_105_port, IN4 => n4995, Q => n1944);
   U1944 : AO22X1 port map( IN1 => n5025, IN2 => RAMDIN1(106), IN3 => 
                           RAM_1_106_port, IN4 => n4995, Q => n1945);
   U1945 : AO22X1 port map( IN1 => n5025, IN2 => RAMDIN1(107), IN3 => 
                           RAM_1_107_port, IN4 => n4995, Q => n1946);
   U1946 : AO22X1 port map( IN1 => n5025, IN2 => RAMDIN1(108), IN3 => 
                           RAM_1_108_port, IN4 => n4995, Q => n1947);
   U1947 : AO22X1 port map( IN1 => n5026, IN2 => RAMDIN1(109), IN3 => 
                           RAM_1_109_port, IN4 => n4995, Q => n1948);
   U1948 : AO22X1 port map( IN1 => RAMDIN1(110), IN2 => n5026, IN3 => 
                           RAM_1_110_port, IN4 => n4995, Q => n1949);
   U1949 : AO22X1 port map( IN1 => n5026, IN2 => RAMDIN1(111), IN3 => 
                           RAM_1_111_port, IN4 => n4995, Q => n1950);
   U1950 : AO22X1 port map( IN1 => RAMDIN1(112), IN2 => n5026, IN3 => 
                           RAM_1_112_port, IN4 => n4995, Q => n1951);
   U1951 : AO22X1 port map( IN1 => n5026, IN2 => RAMDIN1(113), IN3 => 
                           RAM_1_113_port, IN4 => n4995, Q => n1952);
   U1952 : AO22X1 port map( IN1 => n5027, IN2 => RAMDIN1(114), IN3 => 
                           RAM_1_114_port, IN4 => n4995, Q => n1953);
   U1953 : AO22X1 port map( IN1 => RAMDIN1(115), IN2 => n5027, IN3 => 
                           RAM_1_115_port, IN4 => n4995, Q => n1954);
   U1954 : AO22X1 port map( IN1 => n5027, IN2 => RAMDIN1(116), IN3 => 
                           RAM_1_116_port, IN4 => n4994, Q => n1955);
   U1955 : AO22X1 port map( IN1 => n5027, IN2 => RAMDIN1(117), IN3 => 
                           RAM_1_117_port, IN4 => n4994, Q => n1956);
   U1956 : AO22X1 port map( IN1 => n5027, IN2 => RAMDIN1(118), IN3 => 
                           RAM_1_118_port, IN4 => n4994, Q => n1957);
   U1957 : AO22X1 port map( IN1 => n5028, IN2 => RAMDIN1(119), IN3 => 
                           RAM_1_119_port, IN4 => n4994, Q => n1958);
   U1958 : AO22X1 port map( IN1 => n5028, IN2 => RAMDIN1(120), IN3 => 
                           RAM_1_120_port, IN4 => n4994, Q => n1959);
   U1959 : AO22X1 port map( IN1 => n5028, IN2 => RAMDIN1(121), IN3 => 
                           RAM_1_121_port, IN4 => n4994, Q => n1960);
   U1960 : AO22X1 port map( IN1 => n5028, IN2 => RAMDIN1(122), IN3 => 
                           RAM_1_122_port, IN4 => n4994, Q => n1961);
   U1961 : AO22X1 port map( IN1 => n5028, IN2 => RAMDIN1(123), IN3 => 
                           RAM_1_123_port, IN4 => n4994, Q => n1962);
   U1962 : AO22X1 port map( IN1 => n5029, IN2 => RAMDIN1(124), IN3 => 
                           RAM_1_124_port, IN4 => n4994, Q => n1963);
   U1963 : AO22X1 port map( IN1 => n5029, IN2 => RAMDIN1(125), IN3 => 
                           RAM_1_125_port, IN4 => n4994, Q => n1964);
   U1964 : AO22X1 port map( IN1 => n5029, IN2 => RAMDIN1(126), IN3 => 
                           RAM_1_126_port, IN4 => n4994, Q => n1965);
   U1965 : AO22X1 port map( IN1 => RAMDIN1(127), IN2 => n5029, IN3 => 
                           RAM_1_127_port, IN4 => n4994, Q => n1966);
   U1967 : AO22X1 port map( IN1 => n4968, IN2 => RAMDIN1(0), IN3 => 
                           RAM_0_0_port, IN4 => n4962, Q => n1967);
   U1968 : AO22X1 port map( IN1 => n4967, IN2 => RAMDIN1(1), IN3 => 
                           RAM_0_1_port, IN4 => n4962, Q => n1968);
   U1969 : AO22X1 port map( IN1 => n4964, IN2 => RAMDIN1(2), IN3 => 
                           RAM_0_2_port, IN4 => n4962, Q => n1969);
   U1970 : AO22X1 port map( IN1 => n4964, IN2 => RAMDIN1(3), IN3 => 
                           RAM_0_3_port, IN4 => n4962, Q => n1970);
   U1971 : AO22X1 port map( IN1 => n4987, IN2 => RAMDIN1(4), IN3 => 
                           RAM_0_4_port, IN4 => n4962, Q => n1971);
   U1972 : AO22X1 port map( IN1 => n4986, IN2 => RAMDIN1(5), IN3 => 
                           RAM_0_5_port, IN4 => n4962, Q => n1972);
   U1973 : AO22X1 port map( IN1 => n4985, IN2 => RAMDIN1(6), IN3 => 
                           RAM_0_6_port, IN4 => n4962, Q => n1973);
   U1974 : AO22X1 port map( IN1 => RAMDIN1(7), IN2 => n4985, IN3 => 
                           RAM_0_7_port, IN4 => n4962, Q => n1974);
   U1975 : AO22X1 port map( IN1 => RAMDIN1(8), IN2 => n4987, IN3 => 
                           RAM_0_8_port, IN4 => n4961, Q => n1975);
   U1976 : AO22X1 port map( IN1 => n4985, IN2 => RAMDIN1(9), IN3 => 
                           RAM_0_9_port, IN4 => n4961, Q => n1976);
   U1977 : AO22X1 port map( IN1 => n4987, IN2 => RAMDIN1(10), IN3 => 
                           RAM_0_10_port, IN4 => n4961, Q => n1977);
   U1978 : AO22X1 port map( IN1 => RAMDIN1(11), IN2 => n4986, IN3 => 
                           RAM_0_11_port, IN4 => n4961, Q => n1978);
   U1979 : AO22X1 port map( IN1 => RAMDIN1(12), IN2 => n4987, IN3 => 
                           RAM_0_12_port, IN4 => n4961, Q => n1979);
   U1980 : AO22X1 port map( IN1 => n4986, IN2 => RAMDIN1(13), IN3 => 
                           RAM_0_13_port, IN4 => n4961, Q => n1980);
   U1981 : AO22X1 port map( IN1 => RAMDIN1(14), IN2 => n4965, IN3 => 
                           RAM_0_14_port, IN4 => n4961, Q => n1981);
   U1982 : AO22X1 port map( IN1 => n4965, IN2 => RAMDIN1(15), IN3 => 
                           RAM_0_15_port, IN4 => n4961, Q => n1982);
   U1983 : AO22X1 port map( IN1 => RAMDIN1(16), IN2 => n4965, IN3 => 
                           RAM_0_16_port, IN4 => n4961, Q => n1983);
   U1984 : AO22X1 port map( IN1 => n4965, IN2 => RAMDIN1(17), IN3 => 
                           RAM_0_17_port, IN4 => n4961, Q => n1984);
   U1985 : AO22X1 port map( IN1 => RAMDIN1(18), IN2 => n4965, IN3 => 
                           RAM_0_18_port, IN4 => n4961, Q => n1985);
   U1986 : AO22X1 port map( IN1 => n4966, IN2 => RAMDIN1(19), IN3 => 
                           RAM_0_19_port, IN4 => n4961, Q => n1986);
   U1987 : AO22X1 port map( IN1 => RAMDIN1(20), IN2 => n4966, IN3 => 
                           RAM_0_20_port, IN4 => n4960, Q => n1987);
   U1988 : AO22X1 port map( IN1 => n4966, IN2 => RAMDIN1(21), IN3 => 
                           RAM_0_21_port, IN4 => n4960, Q => n1988);
   U1989 : AO22X1 port map( IN1 => n4966, IN2 => n2103, IN3 => RAM_0_22_port, 
                           IN4 => n4960, Q => n1989);
   U1990 : AO22X1 port map( IN1 => n4966, IN2 => RAMDIN1(23), IN3 => 
                           RAM_0_23_port, IN4 => n4960, Q => n1990);
   U1991 : AO22X1 port map( IN1 => n4967, IN2 => n2105, IN3 => RAM_0_24_port, 
                           IN4 => n4960, Q => n1991);
   U1992 : AO22X1 port map( IN1 => n4967, IN2 => RAMDIN1(25), IN3 => 
                           RAM_0_25_port, IN4 => n4960, Q => n1992);
   U1993 : AO22X1 port map( IN1 => n4967, IN2 => RAMDIN1(26), IN3 => 
                           RAM_0_26_port, IN4 => n4960, Q => n1993);
   U1994 : AO22X1 port map( IN1 => n4967, IN2 => RAMDIN1(27), IN3 => 
                           RAM_0_27_port, IN4 => n4960, Q => n1994);
   U1995 : AO22X1 port map( IN1 => RAMDIN1(28), IN2 => n4967, IN3 => 
                           RAM_0_28_port, IN4 => n4960, Q => n1995);
   U1996 : AO22X1 port map( IN1 => n4968, IN2 => RAMDIN1(29), IN3 => 
                           RAM_0_29_port, IN4 => n4960, Q => n1996);
   U1997 : AO22X1 port map( IN1 => n4968, IN2 => RAMDIN1(30), IN3 => 
                           RAM_0_30_port, IN4 => n4960, Q => n1997);
   U1998 : AO22X1 port map( IN1 => n4968, IN2 => RAMDIN1(31), IN3 => 
                           RAM_0_31_port, IN4 => n4960, Q => n1998);
   U1999 : AO22X1 port map( IN1 => n4968, IN2 => RAMDIN1(32), IN3 => 
                           RAM_0_32_port, IN4 => n4959, Q => n1999);
   U2000 : AO22X1 port map( IN1 => n4968, IN2 => RAMDIN1(33), IN3 => 
                           RAM_0_33_port, IN4 => n4959, Q => n2000);
   U2001 : AO22X1 port map( IN1 => RAMDIN1(34), IN2 => n4969, IN3 => 
                           RAM_0_34_port, IN4 => n4959, Q => n2001);
   U2002 : AO22X1 port map( IN1 => n4969, IN2 => RAMDIN1(35), IN3 => 
                           RAM_0_35_port, IN4 => n4959, Q => n2002);
   U2003 : AO22X1 port map( IN1 => n4969, IN2 => RAMDIN1(36), IN3 => 
                           RAM_0_36_port, IN4 => n4959, Q => n2003);
   U2005 : AO22X1 port map( IN1 => n4969, IN2 => RAMDIN1(38), IN3 => 
                           RAM_0_38_port, IN4 => n4959, Q => n2005);
   U2006 : AO22X1 port map( IN1 => n4970, IN2 => RAMDIN1(39), IN3 => 
                           RAM_0_39_port, IN4 => n4959, Q => n2006);
   U2007 : AO22X1 port map( IN1 => RAMDIN1(40), IN2 => n4970, IN3 => 
                           RAM_0_40_port, IN4 => n4959, Q => n2007);
   U2008 : AO22X1 port map( IN1 => n4970, IN2 => n2104, IN3 => RAM_0_41_port, 
                           IN4 => n4959, Q => n2008);
   U2009 : AO22X1 port map( IN1 => n4970, IN2 => RAMDIN1(42), IN3 => 
                           RAM_0_42_port, IN4 => n4959, Q => n2009);
   U2010 : AO22X1 port map( IN1 => n4970, IN2 => n2101, IN3 => RAM_0_43_port, 
                           IN4 => n4959, Q => n2010);
   U2011 : AO22X1 port map( IN1 => n4971, IN2 => RAMDIN1(44), IN3 => 
                           RAM_0_44_port, IN4 => n4958, Q => n2011);
   U2012 : AO22X1 port map( IN1 => n4971, IN2 => RAMDIN1(45), IN3 => 
                           RAM_0_45_port, IN4 => n4958, Q => n2012);
   U2013 : AO22X1 port map( IN1 => RAMDIN1(46), IN2 => n4971, IN3 => 
                           RAM_0_46_port, IN4 => n4958, Q => n2013);
   U2014 : AO22X1 port map( IN1 => RAMDIN1(47), IN2 => n4971, IN3 => 
                           RAM_0_47_port, IN4 => n4958, Q => n2014);
   U2015 : AO22X1 port map( IN1 => n4971, IN2 => n2557, IN3 => RAM_0_48_port, 
                           IN4 => n4958, Q => n2015);
   U2016 : AO22X1 port map( IN1 => RAMDIN1(49), IN2 => n4972, IN3 => 
                           RAM_0_49_port, IN4 => n4958, Q => n2016);
   U2017 : AO22X1 port map( IN1 => n4972, IN2 => RAMDIN1(50), IN3 => 
                           RAM_0_50_port, IN4 => n4958, Q => n2017);
   U2018 : AO22X1 port map( IN1 => n4972, IN2 => RAMDIN1(51), IN3 => 
                           RAM_0_51_port, IN4 => n4958, Q => n2018);
   U2019 : AO22X1 port map( IN1 => n4972, IN2 => n2556, IN3 => RAM_0_52_port, 
                           IN4 => n4958, Q => n2019);
   U2020 : AO22X1 port map( IN1 => n4972, IN2 => RAMDIN1(53), IN3 => 
                           RAM_0_53_port, IN4 => n4958, Q => n2020);
   U2021 : AO22X1 port map( IN1 => n4973, IN2 => RAMDIN1(54), IN3 => 
                           RAM_0_54_port, IN4 => n4958, Q => n2021);
   U2022 : AO22X1 port map( IN1 => n4973, IN2 => RAMDIN1(55), IN3 => 
                           RAM_0_55_port, IN4 => n4958, Q => n2022);
   U2023 : AO22X1 port map( IN1 => n4973, IN2 => RAMDIN1(56), IN3 => 
                           RAM_0_56_port, IN4 => n4957, Q => n2023);
   U2024 : AO22X1 port map( IN1 => n4973, IN2 => RAMDIN1(57), IN3 => 
                           RAM_0_57_port, IN4 => n4957, Q => n2024);
   U2025 : AO22X1 port map( IN1 => n4973, IN2 => RAMDIN1(58), IN3 => 
                           RAM_0_58_port, IN4 => n4957, Q => n2025);
   U2026 : AO22X1 port map( IN1 => n4974, IN2 => RAMDIN1(59), IN3 => 
                           RAM_0_59_port, IN4 => n4957, Q => n2026);
   U2027 : AO22X1 port map( IN1 => n4974, IN2 => RAMDIN1(60), IN3 => 
                           RAM_0_60_port, IN4 => n4957, Q => n2027);
   U2028 : AO22X1 port map( IN1 => n4974, IN2 => RAMDIN1(61), IN3 => 
                           RAM_0_61_port, IN4 => n4957, Q => n2028);
   U2029 : AO22X1 port map( IN1 => n4974, IN2 => RAMDIN1(62), IN3 => 
                           RAM_0_62_port, IN4 => n4957, Q => n2029);
   U2030 : AO22X1 port map( IN1 => n4974, IN2 => RAMDIN1(63), IN3 => 
                           RAM_0_63_port, IN4 => n4957, Q => n2030);
   U2031 : AO22X1 port map( IN1 => n4975, IN2 => RAMDIN1(64), IN3 => 
                           RAM_0_64_port, IN4 => n4957, Q => n2031);
   U2032 : AO22X1 port map( IN1 => n4975, IN2 => RAMDIN1(65), IN3 => 
                           RAM_0_65_port, IN4 => n4957, Q => n2032);
   U2033 : AO22X1 port map( IN1 => n4975, IN2 => RAMDIN1(66), IN3 => 
                           RAM_0_66_port, IN4 => n4957, Q => n2033);
   U2034 : AO22X1 port map( IN1 => n4975, IN2 => RAMDIN1(67), IN3 => 
                           RAM_0_67_port, IN4 => n4957, Q => n2034);
   U2035 : AO22X1 port map( IN1 => RAMDIN1(68), IN2 => n4975, IN3 => 
                           RAM_0_68_port, IN4 => n4956, Q => n2035);
   U2036 : AO22X1 port map( IN1 => n4976, IN2 => RAMDIN1(69), IN3 => 
                           RAM_0_69_port, IN4 => n4956, Q => n2036);
   U2037 : AO22X1 port map( IN1 => n4976, IN2 => RAMDIN1(70), IN3 => 
                           RAM_0_70_port, IN4 => n4956, Q => n2037);
   U2038 : AO22X1 port map( IN1 => n4976, IN2 => RAMDIN1(71), IN3 => 
                           RAM_0_71_port, IN4 => n4956, Q => n2038);
   U2039 : AO22X1 port map( IN1 => RAMDIN1(72), IN2 => n4976, IN3 => 
                           RAM_0_72_port, IN4 => n4956, Q => n2039);
   U2040 : AO22X1 port map( IN1 => n4976, IN2 => RAMDIN1(73), IN3 => 
                           RAM_0_73_port, IN4 => n4956, Q => n2040);
   U2041 : AO22X1 port map( IN1 => n4977, IN2 => RAMDIN1(74), IN3 => 
                           RAM_0_74_port, IN4 => n4956, Q => n2041);
   U2042 : AO22X1 port map( IN1 => n4977, IN2 => RAMDIN1(75), IN3 => 
                           RAM_0_75_port, IN4 => n4956, Q => n2042);
   U2043 : AO22X1 port map( IN1 => n4977, IN2 => RAMDIN1(76), IN3 => 
                           RAM_0_76_port, IN4 => n4956, Q => n2043);
   U2044 : AO22X1 port map( IN1 => n4977, IN2 => RAMDIN1(77), IN3 => 
                           RAM_0_77_port, IN4 => n4956, Q => n2044);
   U2045 : AO22X1 port map( IN1 => RAMDIN1(78), IN2 => n4977, IN3 => 
                           RAM_0_78_port, IN4 => n4956, Q => n2045);
   U2046 : AO22X1 port map( IN1 => n4978, IN2 => RAMDIN1(79), IN3 => 
                           RAM_0_79_port, IN4 => n4956, Q => n2046);
   U2047 : AO22X1 port map( IN1 => RAMDIN1(80), IN2 => n4978, IN3 => 
                           RAM_0_80_port, IN4 => n4955, Q => n2047);
   U2048 : AO22X1 port map( IN1 => n4978, IN2 => RAMDIN1(81), IN3 => 
                           RAM_0_81_port, IN4 => n4955, Q => n2048);
   U2049 : AO22X1 port map( IN1 => n4978, IN2 => RAMDIN1(82), IN3 => 
                           RAM_0_82_port, IN4 => n4955, Q => n2049);
   U2050 : AO22X1 port map( IN1 => n4978, IN2 => RAMDIN1(83), IN3 => 
                           RAM_0_83_port, IN4 => n4955, Q => n2050);
   U2051 : AO22X1 port map( IN1 => RAMDIN1(84), IN2 => n4979, IN3 => 
                           RAM_0_84_port, IN4 => n4955, Q => n2051);
   U2052 : AO22X1 port map( IN1 => n4979, IN2 => RAMDIN1(85), IN3 => 
                           RAM_0_85_port, IN4 => n4955, Q => n2052);
   U2053 : AO22X1 port map( IN1 => n4979, IN2 => RAMDIN1(86), IN3 => 
                           RAM_0_86_port, IN4 => n4955, Q => n2053);
   U2054 : AO22X1 port map( IN1 => n4979, IN2 => RAMDIN1(87), IN3 => 
                           RAM_0_87_port, IN4 => n4955, Q => n2054);
   U2055 : AO22X1 port map( IN1 => RAMDIN1(88), IN2 => n4979, IN3 => 
                           RAM_0_88_port, IN4 => n4955, Q => n2055);
   U2056 : AO22X1 port map( IN1 => n4980, IN2 => RAMDIN1(89), IN3 => 
                           RAM_0_89_port, IN4 => n4955, Q => n2056);
   U2057 : AO22X1 port map( IN1 => n4980, IN2 => RAMDIN1(90), IN3 => 
                           RAM_0_90_port, IN4 => n4955, Q => n2057);
   U2058 : AO22X1 port map( IN1 => n4980, IN2 => RAMDIN1(91), IN3 => 
                           RAM_0_91_port, IN4 => n4955, Q => n2058);
   U2059 : AO22X1 port map( IN1 => RAMDIN1(92), IN2 => n4980, IN3 => 
                           RAM_0_92_port, IN4 => n4954, Q => n2059);
   U2060 : AO22X1 port map( IN1 => n4980, IN2 => RAMDIN1(93), IN3 => 
                           RAM_0_93_port, IN4 => n4954, Q => n2060);
   U2061 : AO22X1 port map( IN1 => n4981, IN2 => RAMDIN1(94), IN3 => 
                           RAM_0_94_port, IN4 => n4954, Q => n2061);
   U2062 : AO22X1 port map( IN1 => n4981, IN2 => RAMDIN1(95), IN3 => 
                           RAM_0_95_port, IN4 => n4954, Q => n2062);
   U2063 : AO22X1 port map( IN1 => n4981, IN2 => RAMDIN1(96), IN3 => 
                           RAM_0_96_port, IN4 => n4954, Q => n2063);
   U2064 : AO22X1 port map( IN1 => n4981, IN2 => RAMDIN1(97), IN3 => 
                           RAM_0_97_port, IN4 => n4954, Q => n2064);
   U2065 : AO22X1 port map( IN1 => n4981, IN2 => RAMDIN1(98), IN3 => 
                           RAM_0_98_port, IN4 => n4954, Q => n2065);
   U2066 : AO22X1 port map( IN1 => n4982, IN2 => n2102, IN3 => RAM_0_99_port, 
                           IN4 => n4954, Q => n2066);
   U2067 : AO22X1 port map( IN1 => n4982, IN2 => RAMDIN1(100), IN3 => 
                           RAM_0_100_port, IN4 => n4954, Q => n2067);
   U2068 : AO22X1 port map( IN1 => n4982, IN2 => RAMDIN1(101), IN3 => 
                           RAM_0_101_port, IN4 => n4954, Q => n2068);
   U2069 : AO22X1 port map( IN1 => n4982, IN2 => RAMDIN1(102), IN3 => 
                           RAM_0_102_port, IN4 => n4954, Q => n2069);
   U2070 : AO22X1 port map( IN1 => n4982, IN2 => RAMDIN1(103), IN3 => 
                           RAM_0_103_port, IN4 => n4954, Q => n2070);
   U2071 : AO22X1 port map( IN1 => n4983, IN2 => RAMDIN1(104), IN3 => 
                           RAM_0_104_port, IN4 => n4953, Q => n2071);
   U2072 : AO22X1 port map( IN1 => n4983, IN2 => RAMDIN1(105), IN3 => 
                           RAM_0_105_port, IN4 => n4953, Q => n2072);
   U2073 : AO22X1 port map( IN1 => n4983, IN2 => RAMDIN1(106), IN3 => 
                           RAM_0_106_port, IN4 => n4953, Q => n2073);
   U2074 : AO22X1 port map( IN1 => n4983, IN2 => RAMDIN1(107), IN3 => 
                           RAM_0_107_port, IN4 => n4953, Q => n2074);
   U2075 : AO22X1 port map( IN1 => n4983, IN2 => RAMDIN1(108), IN3 => 
                           RAM_0_108_port, IN4 => n4953, Q => n2075);
   U2076 : AO22X1 port map( IN1 => n4984, IN2 => RAMDIN1(109), IN3 => 
                           RAM_0_109_port, IN4 => n4953, Q => n2076);
   U2077 : AO22X1 port map( IN1 => RAMDIN1(110), IN2 => n4984, IN3 => 
                           RAM_0_110_port, IN4 => n4953, Q => n2077);
   U2078 : AO22X1 port map( IN1 => n4984, IN2 => RAMDIN1(111), IN3 => 
                           RAM_0_111_port, IN4 => n4953, Q => n2078);
   U2079 : AO22X1 port map( IN1 => RAMDIN1(112), IN2 => n4984, IN3 => 
                           RAM_0_112_port, IN4 => n4953, Q => n2079);
   U2080 : AO22X1 port map( IN1 => RAMDIN1(113), IN2 => n4984, IN3 => 
                           RAM_0_113_port, IN4 => n4953, Q => n2080);
   U2081 : AO22X1 port map( IN1 => n4985, IN2 => RAMDIN1(114), IN3 => 
                           RAM_0_114_port, IN4 => n4953, Q => n2081);
   U2082 : AO22X1 port map( IN1 => n4985, IN2 => RAMDIN1(115), IN3 => 
                           RAM_0_115_port, IN4 => n4953, Q => n2082);
   U2083 : AO22X1 port map( IN1 => n4985, IN2 => RAMDIN1(116), IN3 => 
                           RAM_0_116_port, IN4 => n4952, Q => n2083);
   U2084 : AO22X1 port map( IN1 => n4985, IN2 => RAMDIN1(117), IN3 => 
                           RAM_0_117_port, IN4 => n4952, Q => n2084);
   U2085 : AO22X1 port map( IN1 => n4985, IN2 => RAMDIN1(118), IN3 => 
                           RAM_0_118_port, IN4 => n4952, Q => n2085);
   U2086 : AO22X1 port map( IN1 => n4986, IN2 => RAMDIN1(119), IN3 => 
                           RAM_0_119_port, IN4 => n4952, Q => n2086);
   U2087 : AO22X1 port map( IN1 => RAMDIN1(120), IN2 => n4986, IN3 => 
                           RAM_0_120_port, IN4 => n4952, Q => n2087);
   U2088 : AO22X1 port map( IN1 => n4986, IN2 => RAMDIN1(121), IN3 => 
                           RAM_0_121_port, IN4 => n4952, Q => n2088);
   U2089 : AO22X1 port map( IN1 => n4986, IN2 => RAMDIN1(122), IN3 => 
                           RAM_0_122_port, IN4 => n4952, Q => n2089);
   U2090 : AO22X1 port map( IN1 => n4986, IN2 => RAMDIN1(123), IN3 => 
                           RAM_0_123_port, IN4 => n4952, Q => n2090);
   U2091 : AO22X1 port map( IN1 => n4987, IN2 => RAMDIN1(124), IN3 => 
                           RAM_0_124_port, IN4 => n4952, Q => n2091);
   U2092 : AO22X1 port map( IN1 => n4987, IN2 => RAMDIN1(125), IN3 => 
                           RAM_0_125_port, IN4 => n4952, Q => n2092);
   U2093 : AO22X1 port map( IN1 => n4987, IN2 => RAMDIN1(126), IN3 => 
                           RAM_0_126_port, IN4 => n4952, Q => n2093);
   U2094 : AO22X1 port map( IN1 => RAMDIN1(127), IN2 => n4987, IN3 => 
                           RAM_0_127_port, IN4 => n4952, Q => n2094);
   U2095 : AND2X1 port map( IN1 => n45, IN2 => n2708, Q => n39);
   U2 : AOI221X1 port map( IN1 => RAM_8_90_port, IN2 => n3426, IN3 => 
                           RAM_9_90_port, IN4 => n3369, IN5 => n3187, QN => 
                           n2266);
   U3 : AND2X4 port map( IN1 => n2828, IN2 => n2819, Q => n3339);
   U4 : NBUFFX2 port map( INP => RAMDIN1(37), Z => n1);
   U5 : NBUFFX2 port map( INP => RAMDIN1(52), Z => n2);
   U6 : AOI221X1 port map( IN1 => RAM_0_97_port, IN2 => n2160, IN3 => 
                           RAM_1_97_port, IN4 => n2492, IN5 => n3217, QN => 
                           n2308);
   U7 : NAND4X0 port map( IN1 => n3, IN2 => n4, IN3 => n5, IN4 => n6, QN => 
                           RAMDOUT1(33));
   U8 : AOI221X1 port map( IN1 => RAM_8_33_port, IN2 => n3421, IN3 => 
                           RAM_9_33_port, IN4 => n3369, IN5 => n2959, QN => n3)
                           ;
   U9 : AOI221X1 port map( IN1 => RAM_12_33_port, IN2 => n2455, IN3 => n3374, 
                           IN4 => RAM_13_33_port, IN5 => n2960, QN => n4);
   U10 : AOI221X1 port map( IN1 => RAM_0_33_port, IN2 => n2170, IN3 => n3382, 
                           IN4 => RAM_1_33_port, IN5 => n2961, QN => n5);
   U11 : AOI221X2 port map( IN1 => RAM_4_33_port, IN2 => n3405, IN3 => 
                           RAM_5_33_port, IN4 => n3401, IN5 => n2962, QN => n6)
                           ;
   U12 : AOI221X1 port map( IN1 => RAM_8_3_port, IN2 => n3415, IN3 => 
                           RAM_9_3_port, IN4 => n3363, IN5 => n2839, QN => 
                           n3414);
   U13 : AOI221X1 port map( IN1 => RAM_0_9_port, IN2 => n2166, IN3 => 
                           RAM_1_9_port, IN4 => n2157, IN5 => n2865, QN => 
                           n2292);
   U14 : AO22X1 port map( IN1 => RAM_15_91_port, IN2 => n3441, IN3 => 
                           RAM_14_91_port, IN4 => n2331, Q => n3192);
   U15 : AOI221X1 port map( IN1 => RAM_0_101_port, IN2 => n2170, IN3 => 
                           RAM_1_101_port, IN4 => n3386, IN5 => n3233, QN => 
                           n2736);
   U16 : AOI221X1 port map( IN1 => RAM_0_107_port, IN2 => n2173, IN3 => 
                           RAM_1_107_port, IN4 => n3383, IN5 => n3257, QN => 
                           n2712);
   U17 : AOI221X1 port map( IN1 => RAM_0_45_port, IN2 => n2165, IN3 => 
                           RAM_1_45_port, IN4 => n2157, IN5 => n3009, QN => 
                           n2588);
   U18 : AOI221X1 port map( IN1 => RAM_0_55_port, IN2 => n2168, IN3 => 
                           RAM_1_55_port, IN4 => n3387, IN5 => n3049, QN => 
                           n2234);
   U19 : AO22X1 port map( IN1 => RAM_15_59_port, IN2 => n3443, IN3 => 
                           RAM_14_59_port, IN4 => n2338, Q => n3064);
   U20 : AO22X1 port map( IN1 => RAM_15_82_port, IN2 => n3443, IN3 => 
                           RAM_14_82_port, IN4 => n2334, Q => n3156);
   U21 : AO22X1 port map( IN1 => RAM_15_113_port, IN2 => n3443, IN3 => 
                           RAM_14_113_port, IN4 => n2332, Q => n3284);
   U22 : AO22X1 port map( IN1 => RAM_15_76_port, IN2 => n3443, IN3 => 
                           RAM_14_76_port, IN4 => n2323, Q => n3132);
   U23 : AO22X1 port map( IN1 => RAM_15_71_port, IN2 => n3443, IN3 => 
                           RAM_14_71_port, IN4 => n2338, Q => n3112);
   U24 : AO22X1 port map( IN1 => RAM_15_61_port, IN2 => n3443, IN3 => 
                           RAM_14_61_port, IN4 => n2334, Q => n3072);
   U25 : AO22X1 port map( IN1 => RAM_15_97_port, IN2 => n3443, IN3 => 
                           RAM_14_97_port, IN4 => n2327, Q => n3216);
   U26 : AO22X1 port map( IN1 => RAM_15_35_port, IN2 => n3443, IN3 => 
                           RAM_14_35_port, IN4 => n2335, Q => n2968);
   U27 : AOI221X1 port map( IN1 => RAM_0_23_port, IN2 => n2159, IN3 => 
                           RAM_1_23_port, IN4 => n3386, IN5 => n2921, QN => 
                           n2194);
   U28 : DELLN1X2 port map( INP => n3447, Z => n3443);
   U29 : DELLN1X2 port map( INP => n3447, Z => n3437);
   U30 : DELLN1X2 port map( INP => n3447, Z => n3435);
   U31 : DELLN1X2 port map( INP => n3447, Z => n3438);
   U32 : DELLN1X2 port map( INP => n3447, Z => n3433);
   U33 : DELLN1X2 port map( INP => n3447, Z => n3434);
   U34 : DELLN1X2 port map( INP => n3447, Z => n3432);
   U35 : DELLN1X2 port map( INP => n3447, Z => n3436);
   U36 : AOI221X1 port map( IN1 => RAM_12_51_port, IN2 => n2449, IN3 => 
                           RAM_13_51_port, IN4 => n2490, IN5 => n3032, QN => 
                           n2681);
   U37 : AO22X1 port map( IN1 => RAM_15_51_port, IN2 => n3443, IN3 => 
                           RAM_14_51_port, IN4 => n2320, Q => n3032);
   U38 : AOI221X1 port map( IN1 => RAM_12_126_port, IN2 => n2458, IN3 => 
                           RAM_13_126_port, IN4 => n2490, IN5 => n3336, QN => 
                           n2739);
   U39 : AO22X1 port map( IN1 => RAM_15_110_port, IN2 => n3444, IN3 => 
                           RAM_14_110_port, IN4 => n2324, Q => n3268);
   U40 : NBUFFX2 port map( INP => n2318, Z => n2324);
   U41 : AOI221X1 port map( IN1 => RAM_12_83_port, IN2 => n2447, IN3 => 
                           RAM_13_83_port, IN4 => n2490, IN5 => n3160, QN => 
                           n2255);
   U42 : AND2X2 port map( IN1 => n2819, IN2 => n2826, Q => n3342);
   U99 : AND2X1 port map( IN1 => n2825, IN2 => n2829, Q => n3357);
   U100 : NBUFFX2 port map( INP => n2743, Z => n2136);
   U101 : NBUFFX4 port map( INP => n2742, Z => n2142);
   U227 : INVX0 port map( INP => n16, ZN => n3453);
   U228 : INVX0 port map( INP => n16, ZN => n3451);
   U229 : AND2X4 port map( IN1 => n2825, IN2 => n2823, Q => n3352);
   U230 : AO22X2 port map( IN1 => RAM_3_57_port, IN2 => n2537, IN3 => n2644, 
                           IN4 => RAM_2_57_port, Q => n3057);
   U231 : AOI221X1 port map( IN1 => RAM_8_14_port, IN2 => n3418, IN3 => 
                           RAM_9_14_port, IN4 => n3363, IN5 => n2883, QN => 
                           n2578);
   U232 : AO22X1 port map( IN1 => RAM_15_70_port, IN2 => n3442, IN3 => 
                           RAM_14_70_port, IN4 => n2334, Q => n3108);
   U233 : AO22X1 port map( IN1 => RAM_15_18_port, IN2 => n3442, IN3 => 
                           RAM_14_18_port, IN4 => n2338, Q => n2900);
   U234 : AO22X1 port map( IN1 => RAM_15_27_port, IN2 => n3442, IN3 => 
                           RAM_14_27_port, IN4 => n2332, Q => n2936);
   U235 : AO22X1 port map( IN1 => RAM_15_87_port, IN2 => n3442, IN3 => 
                           RAM_14_87_port, IN4 => n2336, Q => n3176);
   U236 : AO22X1 port map( IN1 => RAM_15_112_port, IN2 => n3442, IN3 => 
                           RAM_14_112_port, IN4 => n2339, Q => n3276);
   U237 : AO22X1 port map( IN1 => RAM_15_14_port, IN2 => n3442, IN3 => 
                           RAM_14_14_port, IN4 => n2332, Q => n2884);
   U238 : AOI221X1 port map( IN1 => RAM_0_83_port, IN2 => n2172, IN3 => 
                           RAM_1_83_port, IN4 => n2121, IN5 => n3161, QN => 
                           n2256);
   U939 : AOI221X1 port map( IN1 => RAM_8_80_port, IN2 => n3421, IN3 => 
                           RAM_9_80_port, IN4 => n3361, IN5 => n3147, QN => 
                           n2471);
   U1068 : AOI221X1 port map( IN1 => RAM_0_66_port, IN2 => n2164, IN3 => 
                           RAM_1_66_port, IN4 => n2121, IN5 => n3093, QN => 
                           n2185);
   U1069 : INVX0 port map( INP => n2619, ZN => n7);
   U1250 : AO22X2 port map( IN1 => RAM_3_118_port, IN2 => n2543, IN3 => 
                           RAM_2_118_port, IN4 => n2639, Q => n3305);
   U1966 : AO22X2 port map( IN1 => RAM_3_56_port, IN2 => n2500, IN3 => 
                           RAM_2_56_port, IN4 => n2641, Q => n3053);
   U2004 : AO22X2 port map( IN1 => RAM_3_30_port, IN2 => n2548, IN3 => 
                           RAM_2_30_port, IN4 => n2632, Q => n2949);
   U2096 : AO22X2 port map( IN1 => RAM_3_6_port, IN2 => n2547, IN3 => 
                           RAM_2_6_port, IN4 => n2099, Q => n2853);
   U2097 : AO22X2 port map( IN1 => RAM_11_46_port, IN2 => n3461, IN3 => 
                           RAM_10_46_port, IN4 => n2664, Q => n3011);
   U2098 : IBUFFX16 port map( INP => RAMADDR1(0), ZN => n2708);
   U2099 : AOI221X1 port map( IN1 => RAM_12_89_port, IN2 => n2448, IN3 => 
                           RAM_13_89_port, IN4 => n3380, IN5 => n3184, QN => 
                           n2251);
   U2100 : AOI221X1 port map( IN1 => RAM_8_46_port, IN2 => n3417, IN3 => 
                           RAM_9_46_port, IN4 => n3360, IN5 => n3011, QN => 
                           n2424);
   U2101 : NAND4X0 port map( IN1 => n8, IN2 => n9, IN3 => n10, IN4 => n11, QN 
                           => RAMDOUT1(57));
   U2102 : AOI221X1 port map( IN1 => RAM_8_57_port, IN2 => n3426, IN3 => 
                           RAM_9_57_port, IN4 => n2493, IN5 => n3055, QN => n8)
                           ;
   U2103 : AOI221X1 port map( IN1 => RAM_12_57_port, IN2 => n2454, IN3 => 
                           RAM_13_57_port, IN4 => n3372, IN5 => n3056, QN => n9
                           );
   U2104 : AOI221X1 port map( IN1 => RAM_4_57_port, IN2 => n3448, IN3 => 
                           RAM_5_57_port, IN4 => n3394, IN5 => n3058, QN => n10
                           );
   U2105 : AOI221X1 port map( IN1 => RAM_0_57_port, IN2 => n2173, IN3 => 
                           RAM_1_57_port, IN4 => n2121, IN5 => n3057, QN => n11
                           );
   U2106 : AOI221X1 port map( IN1 => RAM_0_58_port, IN2 => n2160, IN3 => 
                           RAM_1_58_port, IN4 => n3385, IN5 => n3061, QN => 
                           n2363);
   U2107 : NAND4X0 port map( IN1 => n12, IN2 => n13, IN3 => n14, IN4 => n15, QN
                           => RAMDOUT1(115));
   U2108 : AOI221X1 port map( IN1 => RAM_8_115_port, IN2 => n3424, IN3 => 
                           RAM_9_115_port, IN4 => n2493, IN5 => n3291, QN => 
                           n12);
   U2109 : AOI221X1 port map( IN1 => RAM_12_115_port, IN2 => n2457, IN3 => 
                           n3373, IN4 => RAM_13_115_port, IN5 => n3292, QN => 
                           n13);
   U2110 : AOI221X1 port map( IN1 => RAM_0_115_port, IN2 => n2160, IN3 => 
                           RAM_1_115_port, IN4 => n2121, IN5 => n3293, QN => 
                           n14);
   U2111 : AOI221X1 port map( IN1 => RAM_4_115_port, IN2 => n3448, IN3 => 
                           RAM_5_115_port, IN4 => n2495, IN5 => n3294, QN => 
                           n15);
   U2112 : NAND2X0 port map( IN1 => n2819, IN2 => n2827, QN => n16);
   U2113 : IBUFFX16 port map( INP => n2532, ZN => n2537);
   U2114 : AND2X2 port map( IN1 => n2823, IN2 => n2827, Q => n3349);
   U2115 : AO22X2 port map( IN1 => RAM_3_96_port, IN2 => n2550, IN3 => n7, IN4 
                           => RAM_2_96_port, Q => n3213);
   U2116 : AOI221X1 port map( IN1 => RAM_0_77_port, IN2 => n2173, IN3 => 
                           RAM_1_77_port, IN4 => n3384, IN5 => n3137, QN => 
                           n2296);
   U2117 : AOI221X1 port map( IN1 => RAM_0_89_port, IN2 => n2172, IN3 => 
                           RAM_1_89_port, IN4 => n3389, IN5 => n3185, QN => 
                           n2252);
   U2118 : NAND4X0 port map( IN1 => n17, IN2 => n18, IN3 => n19, IN4 => n20, QN
                           => RAMDOUT1(74));
   U2119 : AOI221X1 port map( IN1 => RAM_8_74_port, IN2 => n3425, IN3 => 
                           RAM_9_74_port, IN4 => n3365, IN5 => n3123, QN => n17
                           );
   U2120 : AOI221X1 port map( IN1 => RAM_12_74_port, IN2 => n2456, IN3 => 
                           RAM_13_74_port, IN4 => n3371, IN5 => n3124, QN => 
                           n18);
   U2121 : AOI221X1 port map( IN1 => RAM_0_74_port, IN2 => n2160, IN3 => 
                           RAM_1_74_port, IN4 => n3388, IN5 => n3125, QN => n19
                           );
   U2122 : AOI221X1 port map( IN1 => RAM_4_74_port, IN2 => n3448, IN3 => 
                           RAM_5_74_port, IN4 => n3401, IN5 => n3126, QN => n20
                           );
   U2123 : INVX0 port map( INP => n3348, ZN => n2620);
   U2124 : NAND4X0 port map( IN1 => n2095, IN2 => n2096, IN3 => n2097, IN4 => 
                           n2098, QN => RAMDOUT1(88));
   U2125 : AOI221X1 port map( IN1 => RAM_8_88_port, IN2 => n3421, IN3 => 
                           RAM_9_88_port, IN4 => n3367, IN5 => n3179, QN => 
                           n2095);
   U2126 : AOI221X1 port map( IN1 => RAM_12_88_port, IN2 => n2459, IN3 => 
                           RAM_13_88_port, IN4 => n3377, IN5 => n3180, QN => 
                           n2096);
   U2127 : AOI221X1 port map( IN1 => RAM_0_88_port, IN2 => n2171, IN3 => 
                           RAM_1_88_port, IN4 => n2492, IN5 => n3181, QN => 
                           n2097);
   U2128 : AOI221X1 port map( IN1 => RAM_4_88_port, IN2 => n3403, IN3 => 
                           RAM_5_88_port, IN4 => n3395, IN5 => n3182, QN => 
                           n2098);
   U2129 : INVX0 port map( INP => n2620, ZN => n2099);
   U2130 : AO22X2 port map( IN1 => RAM_11_40_port, IN2 => n3461, IN3 => n2654, 
                           IN4 => RAM_10_40_port, Q => n2987);
   U2131 : AO22X2 port map( IN1 => RAM_11_51_port, IN2 => n2498, IN3 => 
                           RAM_10_51_port, IN4 => n2662, Q => n3031);
   U2132 : AO22X2 port map( IN1 => RAM_11_97_port, IN2 => n3456, IN3 => 
                           RAM_10_97_port, IN4 => n2655, Q => n3215);
   U2133 : AO22X2 port map( IN1 => RAM_11_89_port, IN2 => n2498, IN3 => 
                           RAM_10_89_port, IN4 => n2655, Q => n3183);
   U2134 : AO22X2 port map( IN1 => RAM_11_95_port, IN2 => n3459, IN3 => 
                           RAM_10_95_port, IN4 => n2652, Q => n3207);
   U2135 : AO22X2 port map( IN1 => RAM_11_21_port, IN2 => n3452, IN3 => 
                           RAM_10_21_port, IN4 => n2480, Q => n2911);
   U2136 : AO22X2 port map( IN1 => RAM_11_24_port, IN2 => n2466, IN3 => 
                           RAM_10_24_port, IN4 => n2659, Q => n2923);
   U2137 : AO22X2 port map( IN1 => RAM_11_31_port, IN2 => n3462, IN3 => n2658, 
                           IN4 => RAM_10_31_port, Q => n2951);
   U2138 : AO22X2 port map( IN1 => RAM_11_99_port, IN2 => n2498, IN3 => 
                           RAM_10_99_port, IN4 => n2658, Q => n3223);
   U2139 : AO22X2 port map( IN1 => RAM_11_30_port, IN2 => n3449, IN3 => n2658, 
                           IN4 => RAM_10_30_port, Q => n2947);
   U2140 : AO22X2 port map( IN1 => RAM_11_107_port, IN2 => n3456, IN3 => 
                           RAM_10_107_port, IN4 => n2667, Q => n3255);
   U2141 : AO22X2 port map( IN1 => RAM_11_101_port, IN2 => n3462, IN3 => n2373,
                           IN4 => RAM_10_101_port, Q => n3231);
   U2142 : AO22X2 port map( IN1 => RAM_11_87_port, IN2 => n3454, IN3 => 
                           RAM_10_87_port, IN4 => n2653, Q => n3175);
   U2143 : AO22X2 port map( IN1 => RAM_11_13_port, IN2 => n3457, IN3 => 
                           RAM_10_13_port, IN4 => n2660, Q => n2879);
   U2144 : AO22X2 port map( IN1 => RAM_11_28_port, IN2 => n3456, IN3 => 
                           RAM_10_28_port, IN4 => n2660, Q => n2939);
   U2145 : AND2X2 port map( IN1 => RAMADDR1(3), IN2 => n2100, Q => n2821);
   U2146 : NBUFFX2 port map( INP => RAMADDR1(2), Z => n2100);
   U2147 : AND2X1 port map( IN1 => n2826, IN2 => n2202, Q => n3356);
   U2148 : AND2X4 port map( IN1 => n2826, IN2 => n2821, Q => n3346);
   U2149 : IBUFFX16 port map( INP => n16, ZN => n3459);
   U2150 : IBUFFX16 port map( INP => n16, ZN => n3454);
   U2151 : AO22X2 port map( IN1 => RAM_11_55_port, IN2 => n3456, IN3 => n2662, 
                           IN4 => RAM_10_55_port, Q => n3047);
   U2152 : AO22X2 port map( IN1 => RAM_11_74_port, IN2 => n3456, IN3 => n2657, 
                           IN4 => RAM_10_74_port, Q => n3123);
   U2153 : AO22X2 port map( IN1 => RAM_11_57_port, IN2 => n3457, IN3 => 
                           RAM_10_57_port, IN4 => n2651, Q => n3055);
   U2154 : NBUFFX2 port map( INP => n3352, Z => n2173);
   U2155 : NBUFFX2 port map( INP => n3352, Z => n2160);
   U2156 : NBUFFX2 port map( INP => n3347, Z => n2454);
   U2157 : NBUFFX2 port map( INP => n3347, Z => n2460);
   U2158 : AO22X1 port map( IN1 => RAM_7_20_port, IN2 => n2527, IN3 => 
                           RAM_6_20_port, IN4 => n2148, Q => n2910);
   U2159 : AO22X1 port map( IN1 => RAM_7_65_port, IN2 => n2340, IN3 => 
                           RAM_6_65_port, IN4 => n2147, Q => n3090);
   U2160 : AO22X1 port map( IN1 => RAM_7_24_port, IN2 => n2340, IN3 => 
                           RAM_6_24_port, IN4 => n2139, Q => n2926);
   U2161 : AO22X1 port map( IN1 => RAM_7_99_port, IN2 => n2517, IN3 => 
                           RAM_6_99_port, IN4 => n2137, Q => n3226);
   U2162 : AO22X1 port map( IN1 => RAM_7_5_port, IN2 => n2526, IN3 => 
                           RAM_6_5_port, IN4 => n2152, Q => n2850);
   U2163 : AO22X1 port map( IN1 => RAM_7_33_port, IN2 => n2526, IN3 => 
                           RAM_6_33_port, IN4 => n2152, Q => n2962);
   U2164 : AO22X1 port map( IN1 => RAM_7_107_port, IN2 => n2529, IN3 => 
                           RAM_6_107_port, IN4 => n2152, Q => n3258);
   U2165 : AO22X1 port map( IN1 => RAM_7_113_port, IN2 => n2524, IN3 => 
                           RAM_6_113_port, IN4 => n2151, Q => n3286);
   U2166 : AO22X1 port map( IN1 => RAM_7_120_port, IN2 => n2526, IN3 => 
                           RAM_6_120_port, IN4 => n2135, Q => n3314);
   U2167 : AO22X1 port map( IN1 => RAM_7_125_port, IN2 => n2516, IN3 => 
                           RAM_6_125_port, IN4 => n2147, Q => n3334);
   U2168 : OR4X1 port map( IN1 => n3282, IN2 => n3281, IN3 => n3280, IN4 => 
                           n3279, Q => RAMDOUT1(112));
   U2169 : AO22X2 port map( IN1 => n4969, IN2 => n2559, IN3 => RAM_0_37_port, 
                           IN4 => n4959, Q => n2004);
   U2170 : NBUFFX2 port map( INP => RAMDIN1(43), Z => n2101);
   U2171 : NBUFFX2 port map( INP => RAMDIN1(99), Z => n2102);
   U2172 : NBUFFX2 port map( INP => RAMDIN1(22), Z => n2103);
   U2173 : AOI221X1 port map( IN1 => RAM_0_99_port, IN2 => n2169, IN3 => 
                           RAM_1_99_port, IN4 => n2491, IN5 => n3225, QN => 
                           n2217);
   U2174 : NBUFFX2 port map( INP => RAMDIN1(41), Z => n2104);
   U2175 : AO22X2 port map( IN1 => n5223, IN2 => n2556, IN3 => RAM_6_52_port, 
                           IN4 => n5209, Q => n1251);
   U2176 : NBUFFX2 port map( INP => RAMDIN1(24), Z => n2105);
   U2177 : NBUFFX2 port map( INP => RAMDIN1(24), Z => n2106);
   U2178 : AOI221X1 port map( IN1 => RAM_0_7_port, IN2 => n2173, IN3 => 
                           RAM_1_7_port, IN4 => n3386, IN5 => n2857, QN => 
                           n2316);
   U2179 : AO22X2 port map( IN1 => RAM_3_4_port, IN2 => n2399, IN3 => 
                           RAM_2_4_port, IN4 => n2626, Q => n2845);
   U2180 : AO22X2 port map( IN1 => RAM_3_114_port, IN2 => n2542, IN3 => 
                           RAM_2_114_port, IN4 => n2626, Q => n3289);
   U2181 : AO22X2 port map( IN1 => RAM_3_39_port, IN2 => n2551, IN3 => 
                           RAM_2_39_port, IN4 => n2627, Q => n2985);
   U2182 : AO22X2 port map( IN1 => RAM_11_58_port, IN2 => n3457, IN3 => 
                           RAM_10_58_port, IN4 => n2653, Q => n3059);
   U2183 : AOI221X1 port map( IN1 => RAM_8_87_port, IN2 => n3416, IN3 => 
                           RAM_9_87_port, IN4 => n3370, IN5 => n3175, QN => 
                           n2432);
   U2184 : AOI221X1 port map( IN1 => RAM_0_4_port, IN2 => n2171, IN3 => 
                           RAM_1_4_port, IN4 => n3384, IN5 => n2845, QN => 
                           n2592);
   U2185 : AOI221X1 port map( IN1 => RAM_0_79_port, IN2 => n2170, IN3 => 
                           RAM_1_79_port, IN4 => n3386, IN5 => n3145, QN => 
                           n2674);
   U2186 : AO22X2 port map( IN1 => RAM_11_49_port, IN2 => n2504, IN3 => n2666, 
                           IN4 => RAM_10_49_port, Q => n3023);
   U2187 : AO22X2 port map( IN1 => RAM_11_116_port, IN2 => n2504, IN3 => n2666,
                           IN4 => RAM_10_116_port, Q => n3295);
   U2188 : AOI221X1 port map( IN1 => RAM_0_53_port, IN2 => n2165, IN3 => 
                           RAM_1_53_port, IN4 => n2491, IN5 => n3041, QN => 
                           n2670);
   U2189 : AO22X2 port map( IN1 => RAM_3_9_port, IN2 => n2546, IN3 => n2631, 
                           IN4 => RAM_2_9_port, Q => n2865);
   U2190 : AO22X2 port map( IN1 => RAM_3_19_port, IN2 => n2554, IN3 => 
                           RAM_2_19_port, IN4 => n2636, Q => n2905);
   U2191 : AO22X2 port map( IN1 => RAM_3_70_port, IN2 => n2470, IN3 => 
                           RAM_2_70_port, IN4 => n2629, Q => n3109);
   U2192 : AO22X2 port map( IN1 => RAM_11_44_port, IN2 => n3459, IN3 => n2191, 
                           IN4 => RAM_10_44_port, Q => n3003);
   U2193 : AO22X2 port map( IN1 => RAM_11_110_port, IN2 => n3452, IN3 => n2191,
                           IN4 => RAM_10_110_port, Q => n3267);
   U2194 : AO22X2 port map( IN1 => RAM_11_105_port, IN2 => n3452, IN3 => n2191,
                           IN4 => RAM_10_105_port, Q => n3247);
   U2195 : AND2X2 port map( IN1 => RAMADDR1(3), IN2 => n3358, Q => n2819);
   U2196 : AO22X2 port map( IN1 => RAM_11_82_port, IN2 => n3452, IN3 => 
                           RAM_10_82_port, IN4 => n2663, Q => n3155);
   U2197 : AO22X2 port map( IN1 => RAM_11_10_port, IN2 => n2466, IN3 => n2663, 
                           IN4 => RAM_10_10_port, Q => n2867);
   U2198 : AND2X2 port map( IN1 => n2819, IN2 => n2827, Q => n3340);
   U2199 : AO22X2 port map( IN1 => RAM_3_105_port, IN2 => n2541, IN3 => n7, IN4
                           => RAM_2_105_port, Q => n3249);
   U2200 : AO22X2 port map( IN1 => RAM_3_115_port, IN2 => n2500, IN3 => 
                           RAM_2_115_port, IN4 => n2633, Q => n3293);
   U2201 : AOI221X1 port map( IN1 => RAM_8_110_port, IN2 => n3417, IN3 => 
                           RAM_9_110_port, IN4 => n3363, IN5 => n3267, QN => 
                           n2117);
   U2202 : NAND4X0 port map( IN1 => n2107, IN2 => n2108, IN3 => n2109, IN4 => 
                           n2110, QN => RAMDOUT1(95));
   U2203 : AOI221X1 port map( IN1 => RAM_8_95_port, IN2 => n3422, IN3 => 
                           RAM_9_95_port, IN4 => n3361, IN5 => n3207, QN => 
                           n2107);
   U2204 : AOI221X1 port map( IN1 => RAM_12_95_port, IN2 => n2456, IN3 => n3380
                           , IN4 => RAM_13_95_port, IN5 => n3208, QN => n2108);
   U2205 : AOI221X1 port map( IN1 => RAM_0_95_port, IN2 => n2158, IN3 => 
                           RAM_1_95_port, IN4 => n3387, IN5 => n3209, QN => 
                           n2109);
   U2206 : AOI221X1 port map( IN1 => RAM_4_95_port, IN2 => n3409, IN3 => 
                           RAM_5_95_port, IN4 => n2494, IN5 => n3210, QN => 
                           n2110);
   U2207 : AOI221X1 port map( IN1 => RAM_0_38_port, IN2 => n2171, IN3 => 
                           RAM_1_38_port, IN4 => n3388, IN5 => n2981, QN => 
                           n2584);
   U2208 : AOI221X1 port map( IN1 => RAM_0_10_port, IN2 => n2171, IN3 => 
                           RAM_1_10_port, IN4 => n2492, IN5 => n2869, QN => 
                           n2300);
   U2209 : AOI221X1 port map( IN1 => RAM_8_82_port, IN2 => n3426, IN3 => 
                           RAM_9_82_port, IN4 => n3366, IN5 => n3155, QN => 
                           n2428);
   U2210 : AOI221X1 port map( IN1 => RAM_0_26_port, IN2 => n2159, IN3 => 
                           RAM_1_26_port, IN4 => n3383, IN5 => n2933, QN => 
                           n2759);
   U2211 : AO22X1 port map( IN1 => RAM_7_121_port, IN2 => n2468, IN3 => 
                           RAM_6_121_port, IN4 => n2132, Q => n3318);
   U2212 : AO22X1 port map( IN1 => RAM_7_57_port, IN2 => n2468, IN3 => 
                           RAM_6_57_port, IN4 => n2138, Q => n3058);
   U2213 : AND2X1 port map( IN1 => n2829, IN2 => n2827, Q => n3354);
   U2214 : AO22X2 port map( IN1 => RAM_11_19_port, IN2 => n3451, IN3 => 
                           RAM_10_19_port, IN4 => n2651, Q => n2903);
   U2215 : AOI221X2 port map( IN1 => RAM_8_59_port, IN2 => n3424, IN3 => 
                           RAM_9_59_port, IN4 => n3368, IN5 => n3063, QN => 
                           n2700);
   U2216 : AOI221X2 port map( IN1 => RAM_8_94_port, IN2 => n3419, IN3 => 
                           RAM_9_94_port, IN4 => n3370, IN5 => n3203, QN => 
                           n2610);
   U2217 : AOI221X2 port map( IN1 => RAM_8_97_port, IN2 => n3422, IN3 => 
                           RAM_9_97_port, IN4 => n3362, IN5 => n3215, QN => 
                           n2306);
   U2218 : AOI221X2 port map( IN1 => RAM_12_26_port, IN2 => n2445, IN3 => 
                           RAM_13_26_port, IN4 => n2490, IN5 => n2932, QN => 
                           n2758);
   U2219 : AO221X2 port map( IN1 => RAM_12_112_port, IN2 => n2460, IN3 => 
                           RAM_13_112_port, IN4 => n2490, IN5 => n3276, Q => 
                           n3281);
   U2220 : DELLN1X2 port map( INP => n3357, Z => n3408);
   U2221 : DELLN1X2 port map( INP => n3357, Z => n3402);
   U2222 : DELLN1X2 port map( INP => n3357, Z => n3405);
   U2223 : DELLN1X2 port map( INP => n3357, Z => n3404);
   U2224 : DELLN1X2 port map( INP => n3357, Z => n3403);
   U2225 : DELLN1X2 port map( INP => n3357, Z => n3409);
   U2226 : DELLN1X2 port map( INP => n3357, Z => n3448);
   U2227 : AO22X2 port map( IN1 => RAM_3_35_port, IN2 => n2540, IN3 => n2624, 
                           IN4 => RAM_2_35_port, Q => n2969);
   U2228 : AO22X2 port map( IN1 => RAM_3_78_port, IN2 => n2543, IN3 => n2631, 
                           IN4 => RAM_2_78_port, Q => n3141);
   U2229 : AOI221X2 port map( IN1 => RAM_0_68_port, IN2 => n2171, IN3 => 
                           RAM_1_68_port, IN4 => n2491, IN5 => n3101, QN => 
                           n2787);
   U2230 : AOI221X2 port map( IN1 => RAM_0_63_port, IN2 => n2162, IN3 => 
                           RAM_1_63_port, IN4 => n2491, IN5 => n3081, QN => 
                           n2477);
   U2231 : INVX0 port map( INP => n2646, ZN => n2666);
   U2232 : AOI221X2 port map( IN1 => RAM_4_35_port, IN2 => n3403, IN3 => 
                           RAM_5_35_port, IN4 => n3397, IN5 => n2970, QN => 
                           n2360);
   U2233 : AOI221X2 port map( IN1 => RAM_4_111_port, IN2 => n3404, IN3 => 
                           RAM_5_111_port, IN4 => n3398, IN5 => n3274, QN => 
                           n2261);
   U2234 : AOI221X2 port map( IN1 => RAM_4_121_port, IN2 => n3408, IN3 => 
                           RAM_5_121_port, IN4 => n3395, IN5 => n3318, QN => 
                           n2801);
   U2235 : AOI221X1 port map( IN1 => RAM_0_71_port, IN2 => n2159, IN3 => 
                           RAM_1_71_port, IN4 => n3387, IN5 => n3113, QN => 
                           n2130);
   U2236 : INVX0 port map( INP => n2621, ZN => n2111);
   U2237 : INVX0 port map( INP => n2646, ZN => n2663);
   U2238 : INVX0 port map( INP => n2622, ZN => n2638);
   U2239 : AO22X2 port map( IN1 => RAM_11_65_port, IN2 => n3451, IN3 => 
                           RAM_10_65_port, IN4 => n2461, Q => n3087);
   U2240 : AO22X2 port map( IN1 => RAM_11_52_port, IN2 => n3454, IN3 => 
                           RAM_10_52_port, IN4 => n2461, Q => n3035);
   U2241 : AO22X2 port map( IN1 => RAM_11_117_port, IN2 => n3461, IN3 => 
                           RAM_10_117_port, IN4 => n2663, Q => n3299);
   U2242 : AO22X2 port map( IN1 => RAM_11_15_port, IN2 => n3462, IN3 => 
                           RAM_10_15_port, IN4 => n2663, Q => n2887);
   U2243 : AOI221X1 port map( IN1 => RAM_8_56_port, IN2 => n3415, IN3 => 
                           RAM_9_56_port, IN4 => n3367, IN5 => n3051, QN => 
                           n2602);
   U2244 : AOI221X1 port map( IN1 => RAM_8_122_port, IN2 => n3420, IN3 => 
                           RAM_9_122_port, IN4 => n3369, IN5 => n3319, QN => 
                           n2481);
   U2245 : AOI221X1 port map( IN1 => RAM_8_65_port, IN2 => n3420, IN3 => 
                           RAM_9_65_port, IN4 => n3362, IN5 => n3087, QN => 
                           n2386);
   U2246 : AOI221X1 port map( IN1 => RAM_8_52_port, IN2 => n3418, IN3 => 
                           RAM_9_52_port, IN4 => n3368, IN5 => n3035, QN => 
                           n2175);
   U2247 : INVX0 port map( INP => n2622, ZN => n2634);
   U2248 : INVX0 port map( INP => n2649, ZN => n2112);
   U2249 : NAND4X0 port map( IN1 => n2113, IN2 => n2114, IN3 => n2115, IN4 => 
                           n2116, QN => RAMDOUT1(21));
   U2250 : AOI221X1 port map( IN1 => RAM_8_21_port, IN2 => n3417, IN3 => 
                           RAM_9_21_port, IN4 => n3360, IN5 => n2911, QN => 
                           n2113);
   U2251 : AOI221X1 port map( IN1 => RAM_12_21_port, IN2 => n2457, IN3 => n3379
                           , IN4 => RAM_13_21_port, IN5 => n2912, QN => n2114);
   U2252 : AOI221X1 port map( IN1 => RAM_0_21_port, IN2 => n2161, IN3 => 
                           RAM_1_21_port, IN4 => n2491, IN5 => n2913, QN => 
                           n2115);
   U2253 : AOI221X1 port map( IN1 => RAM_4_21_port, IN2 => n3408, IN3 => 
                           RAM_5_21_port, IN4 => n3396, IN5 => n2914, QN => 
                           n2116);
   U2254 : NAND4X0 port map( IN1 => n2117, IN2 => n2118, IN3 => n2120, IN4 => 
                           n2119, QN => RAMDOUT1(110));
   U2255 : AOI221X1 port map( IN1 => RAM_12_110_port, IN2 => n2457, IN3 => 
                           RAM_13_110_port, IN4 => n3376, IN5 => n3268, QN => 
                           n2118);
   U2256 : AOI221X1 port map( IN1 => RAM_0_110_port, IN2 => n2163, IN3 => 
                           RAM_1_110_port, IN4 => n3388, IN5 => n3269, QN => 
                           n2119);
   U2257 : AOI221X2 port map( IN1 => RAM_4_110_port, IN2 => n3404, IN3 => 
                           RAM_5_110_port, IN4 => n3400, IN5 => n3270, QN => 
                           n2120);
   U2258 : AO22X2 port map( IN1 => RAM_3_28_port, IN2 => n2544, IN3 => 
                           RAM_2_28_port, IN4 => n2637, Q => n2941);
   U2259 : AO22X2 port map( IN1 => RAM_3_81_port, IN2 => n2547, IN3 => n2637, 
                           IN4 => RAM_2_81_port, Q => n3153);
   U2260 : AO22X2 port map( IN1 => RAM_3_41_port, IN2 => n2500, IN3 => 
                           RAM_2_41_port, IN4 => n2637, Q => n2993);
   U2261 : AO22X2 port map( IN1 => RAM_3_109_port, IN2 => n2500, IN3 => 
                           RAM_2_109_port, IN4 => n2638, Q => n3265);
   U2262 : AO22X2 port map( IN1 => RAM_3_103_port, IN2 => n2500, IN3 => 
                           RAM_2_103_port, IN4 => n2638, Q => n3241);
   U2263 : AOI221X1 port map( IN1 => RAM_8_69_port, IN2 => n3415, IN3 => 
                           RAM_9_69_port, IN4 => n3369, IN5 => n3103, QN => 
                           n2726);
   U2264 : AOI221X1 port map( IN1 => RAM_8_73_port, IN2 => n3425, IN3 => 
                           RAM_9_73_port, IN4 => n3360, IN5 => n3119, QN => 
                           n2374);
   U2265 : AOI221X1 port map( IN1 => RAM_8_7_port, IN2 => n3419, IN3 => 
                           RAM_9_7_port, IN4 => n3364, IN5 => n2855, QN => 
                           n2314);
   U2266 : AOI221X1 port map( IN1 => RAM_8_106_port, IN2 => n3425, IN3 => 
                           RAM_9_106_port, IN4 => n3365, IN5 => n3251, QN => 
                           n2485);
   U2267 : AOI221X1 port map( IN1 => RAM_8_96_port, IN2 => n3415, IN3 => 
                           RAM_9_96_port, IN4 => n3368, IN5 => n3211, QN => 
                           n2274);
   U2268 : AOI221X1 port map( IN1 => RAM_8_17_port, IN2 => n3416, IN3 => 
                           RAM_9_17_port, IN4 => n3363, IN5 => n2895, QN => 
                           n2416);
   U2269 : AOI221X1 port map( IN1 => RAM_8_37_port, IN2 => n3422, IN3 => 
                           RAM_9_37_port, IN4 => n3370, IN5 => n2975, QN => 
                           n2196);
   U2270 : AOI221X1 port map( IN1 => RAM_8_66_port, IN2 => n3423, IN3 => 
                           RAM_9_66_port, IN4 => n2493, IN5 => n3091, QN => 
                           n2183);
   U2271 : AOI221X1 port map( IN1 => RAM_8_16_port, IN2 => n3419, IN3 => 
                           RAM_9_16_port, IN4 => n3366, IN5 => n2891, QN => 
                           n2404);
   U2272 : AOI221X1 port map( IN1 => RAM_8_20_port, IN2 => n3419, IN3 => 
                           RAM_9_20_port, IN4 => n2493, IN5 => n2907, QN => 
                           n2574);
   U2273 : AO22X2 port map( IN1 => RAM_11_93_port, IN2 => n3459, IN3 => 
                           RAM_10_93_port, IN4 => n2660, Q => n3199);
   U2274 : AOI221X1 port map( IN1 => RAM_8_105_port, IN2 => n3415, IN3 => 
                           RAM_9_105_port, IN4 => n3370, IN5 => n3247, QN => 
                           n2369);
   U2275 : AOI221X1 port map( IN1 => RAM_8_44_port, IN2 => n3419, IN3 => 
                           RAM_9_44_port, IN4 => n3366, IN5 => n3003, QN => 
                           n2207);
   U2276 : AOI221X1 port map( IN1 => RAM_8_38_port, IN2 => n3417, IN3 => 
                           RAM_9_38_port, IN4 => n3361, IN5 => n2979, QN => 
                           n2582);
   U2277 : AOI221X1 port map( IN1 => RAM_8_4_port, IN2 => n3421, IN3 => 
                           RAM_9_4_port, IN4 => n3367, IN5 => n2843, QN => 
                           n2590);
   U2278 : AOI221X1 port map( IN1 => RAM_8_18_port, IN2 => n3420, IN3 => 
                           RAM_9_18_port, IN4 => n3368, IN5 => n2899, QN => 
                           n2408);
   U2279 : AOI221X1 port map( IN1 => RAM_8_12_port, IN2 => n3415, IN3 => 
                           RAM_9_12_port, IN4 => n3364, IN5 => n2875, QN => 
                           n2365);
   U2280 : AOI221X1 port map( IN1 => RAM_8_58_port, IN2 => n3423, IN3 => 
                           RAM_9_58_port, IN4 => n3368, IN5 => n3059, QN => 
                           n2361);
   U2281 : AOI221X1 port map( IN1 => RAM_8_28_port, IN2 => n3415, IN3 => 
                           RAM_9_28_port, IN4 => n3361, IN5 => n2939, QN => 
                           n2440);
   U2282 : AO22X2 port map( IN1 => RAM_11_36_port, IN2 => n3457, IN3 => 
                           RAM_10_36_port, IN4 => n2662, Q => n2971);
   U2283 : AO22X2 port map( IN1 => n3459, IN2 => RAM_11_6_port, IN3 => 
                           RAM_10_6_port, IN4 => n2656, Q => n2851);
   U2284 : AO22X2 port map( IN1 => n3459, IN2 => RAM_11_8_port, IN3 => 
                           RAM_10_8_port, IN4 => n2657, Q => n2859);
   U2285 : AOI221X1 port map( IN1 => RAM_8_78_port, IN2 => n3416, IN3 => 
                           RAM_9_78_port, IN4 => n3361, IN5 => n3139, QN => 
                           n2676);
   U2286 : AOI221X1 port map( IN1 => RAM_8_109_port, IN2 => n3423, IN3 => 
                           RAM_9_109_port, IN4 => n3361, IN5 => n3263, QN => 
                           n2436);
   U2287 : AOI221X1 port map( IN1 => RAM_8_114_port, IN2 => n3424, IN3 => 
                           RAM_9_114_port, IN4 => n3364, IN5 => n3287, QN => 
                           n2594);
   U2288 : AOI221X1 port map( IN1 => RAM_8_40_port, IN2 => n3423, IN3 => 
                           RAM_9_40_port, IN4 => n3364, IN5 => n2987, QN => 
                           n2345);
   U2289 : AOI221X1 port map( IN1 => RAM_8_55_port, IN2 => n3426, IN3 => 
                           RAM_9_55_port, IN4 => n3363, IN5 => n3047, QN => 
                           n2232);
   U2290 : AOI221X1 port map( IN1 => RAM_8_39_port, IN2 => n3425, IN3 => 
                           RAM_9_39_port, IN4 => n3362, IN5 => n2983, QN => 
                           n2570);
   U2291 : AOI221X1 port map( IN1 => RAM_8_36_port, IN2 => n3417, IN3 => 
                           RAM_9_36_port, IN4 => n3366, IN5 => n2971, QN => 
                           n2349);
   U2292 : AOI221X1 port map( IN1 => RAM_4_127_port, IN2 => n3402, IN3 => 
                           RAM_5_127_port, IN4 => n3393, IN5 => n3355, QN => 
                           n2344);
   U2293 : DELLN1X2 port map( INP => n3351, Z => n2121);
   U2294 : NAND4X0 port map( IN1 => n2122, IN2 => n2123, IN3 => n2124, IN4 => 
                           n2125, QN => RAMDOUT1(104));
   U2295 : AOI221X1 port map( IN1 => RAM_8_104_port, IN2 => n3425, IN3 => 
                           RAM_9_104_port, IN4 => n3367, IN5 => n3243, QN => 
                           n2122);
   U2296 : AOI221X1 port map( IN1 => RAM_12_104_port, IN2 => n2453, IN3 => 
                           RAM_13_104_port, IN4 => n3381, IN5 => n3244, QN => 
                           n2123);
   U2297 : AOI221X1 port map( IN1 => RAM_0_104_port, IN2 => n2162, IN3 => 
                           RAM_1_104_port, IN4 => n3389, IN5 => n3245, QN => 
                           n2124);
   U2298 : AOI221X2 port map( IN1 => RAM_4_104_port, IN2 => n3405, IN3 => 
                           RAM_5_104_port, IN4 => n3396, IN5 => n3246, QN => 
                           n2125);
   U2299 : AOI221X1 port map( IN1 => RAM_8_127_port, IN2 => n3421, IN3 => 
                           RAM_9_127_port, IN4 => n3369, IN5 => n3341, QN => 
                           n2341);
   U2300 : IBUFFX16 port map( INP => n2499, ZN => n2504);
   U2301 : NBUFFX2 port map( INP => RAMDIN1(48), Z => n2126);
   U2302 : NBUFFX2 port map( INP => RAMDIN1(48), Z => n2127);
   U2303 : NAND4X0 port map( IN1 => n2128, IN2 => n2129, IN3 => n2130, IN4 => 
                           n2131, QN => RAMDOUT1(71));
   U2304 : AOI221X1 port map( IN1 => RAM_8_71_port, IN2 => n3416, IN3 => 
                           RAM_9_71_port, IN4 => n3368, IN5 => n3111, QN => 
                           n2128);
   U2305 : AOI221X1 port map( IN1 => RAM_12_71_port, IN2 => n2448, IN3 => 
                           RAM_13_71_port, IN4 => n3378, IN5 => n3112, QN => 
                           n2129);
   U2306 : AOI221X2 port map( IN1 => RAM_4_71_port, IN2 => n3448, IN3 => 
                           RAM_5_71_port, IN4 => n3398, IN5 => n3114, QN => 
                           n2131);
   U2307 : AO22X2 port map( IN1 => RAM_11_17_port, IN2 => n3451, IN3 => n2656, 
                           IN4 => RAM_10_17_port, Q => n2895);
   U2308 : AOI221X1 port map( IN1 => RAM_0_30_port, IN2 => n2165, IN3 => 
                           RAM_1_30_port, IN4 => n2121, IN5 => n2949, QN => 
                           n2189);
   U2309 : INVX0 port map( INP => n2645, ZN => n2654);
   U2310 : NBUFFX2 port map( INP => n2743, Z => n2132);
   U2311 : DELLN1X2 port map( INP => n2743, Z => n2133);
   U2312 : NBUFFX2 port map( INP => n2743, Z => n2134);
   U2313 : NBUFFX2 port map( INP => n2743, Z => n2135);
   U2314 : NBUFFX2 port map( INP => n2174, Z => n2137);
   U2315 : NBUFFX2 port map( INP => n2174, Z => n2138);
   U2316 : NBUFFX2 port map( INP => n2174, Z => n2139);
   U2317 : NBUFFX2 port map( INP => n2174, Z => n2140);
   U2318 : NBUFFX2 port map( INP => n2174, Z => n2141);
   U2319 : NBUFFX2 port map( INP => n2742, Z => n2143);
   U2320 : NBUFFX2 port map( INP => n2742, Z => n2144);
   U2321 : NBUFFX2 port map( INP => n2742, Z => n2145);
   U2322 : NBUFFX2 port map( INP => n2742, Z => n2146);
   U2323 : NBUFFX2 port map( INP => n3353, Z => n2147);
   U2324 : NBUFFX2 port map( INP => n3353, Z => n2148);
   U2325 : NBUFFX2 port map( INP => n3353, Z => n2149);
   U2326 : NBUFFX2 port map( INP => n3353, Z => n2150);
   U2327 : NBUFFX2 port map( INP => n3353, Z => n2151);
   U2328 : NBUFFX2 port map( INP => n3353, Z => n2152);
   U2329 : AO22X2 port map( IN1 => RAM_11_3_port, IN2 => n3457, IN3 => n2667, 
                           IN4 => RAM_10_3_port, Q => n2839);
   U2330 : AOI221X1 port map( IN1 => RAM_8_100_port, IN2 => n3419, IN3 => 
                           RAM_9_100_port, IN4 => n3367, IN5 => n3227, QN => 
                           n2155);
   U2331 : INVX0 port map( INP => n2619, ZN => n2644);
   U2332 : AO22X2 port map( IN1 => RAM_11_7_port, IN2 => n3457, IN3 => n2656, 
                           IN4 => RAM_10_7_port, Q => n2855);
   U2333 : AO22X2 port map( IN1 => RAM_11_41_port, IN2 => n3456, IN3 => n2112, 
                           IN4 => RAM_10_41_port, Q => n2991);
   U2334 : NAND4X0 port map( IN1 => n2153, IN2 => n2154, IN3 => n2155, IN4 => 
                           n2156, QN => RAMDOUT1(100));
   U2335 : AOI221X2 port map( IN1 => RAM_0_100_port, IN2 => n2159, IN3 => 
                           RAM_1_100_port, IN4 => n3389, IN5 => n3229, QN => 
                           n2153);
   U2336 : AOI221X1 port map( IN1 => RAM_12_100_port, IN2 => n2458, IN3 => 
                           n3374, IN4 => RAM_13_100_port, IN5 => n3228, QN => 
                           n2154);
   U2337 : AOI221X2 port map( IN1 => RAM_4_100_port, IN2 => n3410, IN3 => 
                           RAM_5_100_port, IN4 => n3392, IN5 => n3230, QN => 
                           n2156);
   U2338 : AO22X2 port map( IN1 => RAM_11_34_port, IN2 => n3459, IN3 => 
                           RAM_10_34_port, IN4 => n2467, Q => n2963);
   U2339 : AO22X2 port map( IN1 => RAM_11_113_port, IN2 => n3451, IN3 => 
                           RAM_10_113_port, IN4 => n2659, Q => n3283);
   U2340 : AO22X2 port map( IN1 => RAM_11_11_port, IN2 => n2231, IN3 => 
                           RAM_10_11_port, IN4 => n2659, Q => n2871);
   U2341 : AO22X2 port map( IN1 => RAM_11_92_port, IN2 => n3452, IN3 => 
                           RAM_10_92_port, IN4 => n2659, Q => n3195);
   U2342 : AO22X2 port map( IN1 => RAM_11_48_port, IN2 => n3451, IN3 => 
                           RAM_10_48_port, IN4 => n2661, Q => n3019);
   U2343 : AOI221X1 port map( IN1 => RAM_8_1_port, IN2 => n3419, IN3 => 
                           RAM_9_1_port, IN4 => n3367, IN5 => n2831, QN => 
                           n2353);
   U2344 : AOI221X1 port map( IN1 => RAM_8_75_port, IN2 => n3423, IN3 => 
                           RAM_9_75_port, IN4 => n3365, IN5 => n3127, QN => 
                           n2244);
   U2345 : AOI221X1 port map( IN1 => RAM_8_85_port, IN2 => n3424, IN3 => 
                           RAM_9_85_port, IN4 => n3360, IN5 => n3167, QN => 
                           n2236);
   U2346 : AOI221X1 port map( IN1 => RAM_8_11_port, IN2 => n3420, IN3 => 
                           RAM_9_11_port, IN4 => n3366, IN5 => n2871, QN => 
                           n2223);
   U2347 : AOI221X1 port map( IN1 => RAM_8_45_port, IN2 => n3418, IN3 => 
                           RAM_9_45_port, IN4 => n3360, IN5 => n3007, QN => 
                           n2586);
   U2348 : AO22X2 port map( IN1 => RAM_3_97_port, IN2 => n2543, IN3 => 
                           RAM_2_97_port, IN4 => n2636, Q => n3217);
   U2349 : AO22X2 port map( IN1 => RAM_3_10_port, IN2 => n2545, IN3 => n2637, 
                           IN4 => RAM_2_10_port, Q => n2869);
   U2350 : DELLN1X2 port map( INP => n3351, Z => n2157);
   U2351 : NBUFFX2 port map( INP => n3352, Z => n2158);
   U2352 : DELLN1X2 port map( INP => n3352, Z => n2159);
   U2353 : DELLN1X2 port map( INP => n3352, Z => n2161);
   U2354 : DELLN1X2 port map( INP => n3352, Z => n2162);
   U2355 : DELLN1X2 port map( INP => n3352, Z => n2163);
   U2356 : DELLN1X2 port map( INP => n3352, Z => n2164);
   U2357 : DELLN1X2 port map( INP => n3352, Z => n2165);
   U2358 : DELLN1X2 port map( INP => n3352, Z => n2166);
   U2359 : DELLN1X2 port map( INP => n3352, Z => n2167);
   U2360 : DELLN1X2 port map( INP => n3352, Z => n2168);
   U2361 : DELLN1X2 port map( INP => n3352, Z => n2169);
   U2362 : DELLN1X2 port map( INP => n3352, Z => n2170);
   U2363 : DELLN1X2 port map( INP => n3352, Z => n2171);
   U2364 : DELLN1X2 port map( INP => n3352, Z => n2172);
   U2365 : AOI221X1 port map( IN1 => RAM_0_84_port, IN2 => n2166, IN3 => 
                           RAM_1_84_port, IN4 => n2491, IN5 => n3165, QN => 
                           n2724);
   U2366 : AND2X4 port map( IN1 => n2797, IN2 => n2202, Q => n2174);
   U2367 : AOI221X1 port map( IN1 => RAM_4_18_port, IN2 => n3405, IN3 => 
                           RAM_5_18_port, IN4 => n3394, IN5 => n2902, QN => 
                           n2411);
   U2368 : NAND4X0 port map( IN1 => n2175, IN2 => n2176, IN3 => n2177, IN4 => 
                           n2178, QN => RAMDOUT1(52));
   U2369 : AOI221X2 port map( IN1 => RAM_12_52_port, IN2 => n2455, IN3 => 
                           RAM_13_52_port, IN4 => n2490, IN5 => n3036, QN => 
                           n2176);
   U2370 : AOI221X1 port map( IN1 => RAM_0_52_port, IN2 => n2173, IN3 => 
                           RAM_1_52_port, IN4 => n3385, IN5 => n3037, QN => 
                           n2177);
   U2371 : AOI221X1 port map( IN1 => RAM_4_52_port, IN2 => n3408, IN3 => 
                           RAM_5_52_port, IN4 => n2494, IN5 => n3038, QN => 
                           n2178);
   U2372 : NAND4X0 port map( IN1 => n2179, IN2 => n2180, IN3 => n2181, IN4 => 
                           n2182, QN => RAMDOUT1(48));
   U2373 : AOI221X1 port map( IN1 => RAM_8_48_port, IN2 => n3422, IN3 => 
                           RAM_9_48_port, IN4 => n3360, IN5 => n3019, QN => 
                           n2179);
   U2374 : AOI221X2 port map( IN1 => RAM_12_48_port, IN2 => n2454, IN3 => 
                           RAM_13_48_port, IN4 => n3380, IN5 => n3020, QN => 
                           n2180);
   U2375 : AOI221X1 port map( IN1 => RAM_0_48_port, IN2 => n2170, IN3 => 
                           RAM_1_48_port, IN4 => n3382, IN5 => n3021, QN => 
                           n2181);
   U2376 : AOI221X2 port map( IN1 => RAM_4_48_port, IN2 => n3406, IN3 => 
                           RAM_5_48_port, IN4 => n3393, IN5 => n3022, QN => 
                           n2182);
   U2377 : AOI221X1 port map( IN1 => RAM_8_119_port, IN2 => n3420, IN3 => 
                           RAM_9_119_port, IN4 => n3362, IN5 => n3307, QN => 
                           n2242);
   U2378 : AOI221X1 port map( IN1 => RAM_4_119_port, IN2 => n3409, IN3 => 
                           RAM_5_119_port, IN4 => n3398, IN5 => n3310, QN => 
                           n2243);
   U2379 : DELLN1X2 port map( INP => n3357, Z => n3406);
   U2380 : AO22X2 port map( IN1 => RAM_3_74_port, IN2 => n2548, IN3 => 
                           RAM_2_74_port, IN4 => n7, Q => n3125);
   U2381 : AO22X2 port map( IN1 => RAM_3_0_port, IN2 => n2549, IN3 => n2629, 
                           IN4 => RAM_2_0_port, Q => n2824);
   U2382 : NAND4X0 port map( IN1 => n2183, IN2 => n2184, IN3 => n2185, IN4 => 
                           n2186, QN => RAMDOUT1(66));
   U2383 : AOI221X1 port map( IN1 => RAM_12_66_port, IN2 => n2459, IN3 => n3379
                           , IN4 => RAM_13_66_port, IN5 => n3092, QN => n2184);
   U2384 : AOI221X2 port map( IN1 => RAM_4_66_port, IN2 => n3402, IN3 => 
                           RAM_5_66_port, IN4 => n3399, IN5 => n3094, QN => 
                           n2186);
   U2385 : AOI221X1 port map( IN1 => RAM_4_124_port, IN2 => n3407, IN3 => 
                           RAM_5_124_port, IN4 => n3399, IN5 => n3330, QN => 
                           n2721);
   U2386 : NAND4X0 port map( IN1 => n2187, IN2 => n2188, IN3 => n2189, IN4 => 
                           n2190, QN => RAMDOUT1(30));
   U2387 : AOI221X2 port map( IN1 => RAM_8_30_port, IN2 => n3416, IN3 => 
                           RAM_9_30_port, IN4 => n3370, IN5 => n2947, QN => 
                           n2187);
   U2388 : AOI221X1 port map( IN1 => RAM_12_30_port, IN2 => n2449, IN3 => n3379
                           , IN4 => RAM_13_30_port, IN5 => n2948, QN => n2188);
   U2389 : AOI221X1 port map( IN1 => RAM_4_30_port, IN2 => n3402, IN3 => 
                           RAM_5_30_port, IN4 => n2494, IN5 => n2950, QN => 
                           n2190);
   U2390 : INVX0 port map( INP => n2618, ZN => n2643);
   U2391 : AO22X2 port map( IN1 => RAM_3_71_port, IN2 => n2553, IN3 => 
                           RAM_2_71_port, IN4 => n2640, Q => n3113);
   U2392 : AO22X2 port map( IN1 => RAM_3_12_port, IN2 => n2548, IN3 => 
                           RAM_2_12_port, IN4 => n7, Q => n2877);
   U2393 : AO22X2 port map( IN1 => RAM_3_47_port, IN2 => n2537, IN3 => 
                           RAM_2_47_port, IN4 => n2627, Q => n3017);
   U2394 : AO22X2 port map( IN1 => RAM_3_51_port, IN2 => n2545, IN3 => 
                           RAM_2_51_port, IN4 => n2643, Q => n3033);
   U2395 : AOI221X1 port map( IN1 => RAM_0_73_port, IN2 => n2161, IN3 => 
                           RAM_1_73_port, IN4 => n3388, IN5 => n3121, QN => 
                           n2376);
   U2396 : AOI221X1 port map( IN1 => RAM_0_94_port, IN2 => n2168, IN3 => 
                           RAM_1_94_port, IN4 => n3382, IN5 => n3205, QN => 
                           n2611);
   U2397 : AOI221X1 port map( IN1 => RAM_0_20_port, IN2 => n2173, IN3 => 
                           RAM_1_20_port, IN4 => n3382, IN5 => n2909, QN => 
                           n2576);
   U2398 : AOI221X1 port map( IN1 => RAM_0_35_port, IN2 => n2163, IN3 => 
                           RAM_1_35_port, IN4 => n3386, IN5 => n2969, QN => 
                           n2359);
   U2399 : AOI221X1 port map( IN1 => RAM_0_105_port, IN2 => n2162, IN3 => 
                           RAM_1_105_port, IN4 => n2121, IN5 => n3249, QN => 
                           n2371);
   U2400 : AOI221X1 port map( IN1 => RAM_0_85_port, IN2 => n2170, IN3 => 
                           RAM_1_85_port, IN4 => n3390, IN5 => n3169, QN => 
                           n2238);
   U2401 : AOI221X1 port map( IN1 => RAM_0_76_port, IN2 => n2167, IN3 => 
                           RAM_1_76_port, IN4 => n3387, IN5 => n3133, QN => 
                           n2716);
   U2402 : AOI221X1 port map( IN1 => RAM_8_118_port, IN2 => n3423, IN3 => 
                           RAM_9_118_port, IN4 => n3362, IN5 => n3303, QN => 
                           n2598);
   U2403 : INVX0 port map( INP => n2647, ZN => n2191);
   U2404 : NAND4X0 port map( IN1 => n2192, IN2 => n2193, IN3 => n2194, IN4 => 
                           n2195, QN => RAMDOUT1(23));
   U2405 : AOI221X1 port map( IN1 => RAM_8_23_port, IN2 => n3421, IN3 => 
                           RAM_9_23_port, IN4 => n3362, IN5 => n2919, QN => 
                           n2192);
   U2406 : AOI221X1 port map( IN1 => RAM_12_23_port, IN2 => n2455, IN3 => n3377
                           , IN4 => RAM_13_23_port, IN5 => n2920, QN => n2193);
   U2407 : AOI221X2 port map( IN1 => RAM_4_23_port, IN2 => n3406, IN3 => 
                           RAM_5_23_port, IN4 => n3401, IN5 => n2922, QN => 
                           n2195);
   U2408 : AOI221X1 port map( IN1 => RAM_8_35_port, IN2 => n3415, IN3 => 
                           RAM_9_35_port, IN4 => n3367, IN5 => n2967, QN => 
                           n2357);
   U2409 : AOI221X1 port map( IN1 => RAM_8_117_port, IN2 => n3425, IN3 => 
                           RAM_9_117_port, IN4 => n3362, IN5 => n3299, QN => 
                           n2262);
   U2410 : AOI221X1 port map( IN1 => RAM_8_15_port, IN2 => n3418, IN3 => 
                           RAM_9_15_port, IN4 => n3369, IN5 => n2887, QN => 
                           n2420);
   U2411 : AOI221X1 port map( IN1 => RAM_8_10_port, IN2 => n3420, IN3 => 
                           RAM_9_10_port, IN4 => n3369, IN5 => n2867, QN => 
                           n2298);
   U2412 : AND2X2 port map( IN1 => n2828, IN2 => n2823, Q => n3348);
   U2413 : DELLN2X2 port map( INP => n3357, Z => n3410);
   U2414 : DELLN1X2 port map( INP => n3357, Z => n3407);
   U2415 : NAND4X0 port map( IN1 => n2196, IN2 => n2197, IN3 => n2198, IN4 => 
                           n2199, QN => RAMDOUT1(37));
   U2416 : AOI221X2 port map( IN1 => RAM_12_37_port, IN2 => n2457, IN3 => 
                           RAM_13_37_port, IN4 => n3372, IN5 => n2976, QN => 
                           n2197);
   U2417 : AOI221X1 port map( IN1 => RAM_0_37_port, IN2 => n2172, IN3 => 
                           RAM_1_37_port, IN4 => n3382, IN5 => n2977, QN => 
                           n2198);
   U2418 : AOI221X2 port map( IN1 => RAM_4_37_port, IN2 => n3403, IN3 => 
                           RAM_5_37_port, IN4 => n2495, IN5 => n2978, QN => 
                           n2199);
   U2419 : NBUFFX2 port map( INP => RAMDIN1(24), Z => n2200);
   U2420 : NBUFFX2 port map( INP => RAMDIN1(24), Z => n2201);
   U2421 : AO22X2 port map( IN1 => RAM_11_70_port, IN2 => n2501, IN3 => n2665, 
                           IN4 => RAM_10_70_port, Q => n3107);
   U2422 : AO22X2 port map( IN1 => RAM_11_64_port, IN2 => n3453, IN3 => 
                           RAM_10_64_port, IN4 => n2666, Q => n3083);
   U2423 : AO22X2 port map( IN1 => RAM_11_108_port, IN2 => n3459, IN3 => 
                           RAM_10_108_port, IN4 => n2667, Q => n3259);
   U2424 : AO22X2 port map( IN1 => RAM_11_43_port, IN2 => n3457, IN3 => 
                           RAM_10_43_port, IN4 => n2656, Q => n2999);
   U2425 : AOI221X1 port map( IN1 => RAM_8_42_port, IN2 => n3426, IN3 => 
                           RAM_9_42_port, IN4 => n3370, IN5 => n2995, QN => 
                           n2562);
   U2426 : AOI221X1 port map( IN1 => RAM_8_60_port, IN2 => n3416, IN3 => 
                           RAM_9_60_port, IN4 => n3363, IN5 => n3067, QN => 
                           n2286);
   U2427 : AOI221X1 port map( IN1 => RAM_8_9_port, IN2 => n3417, IN3 => 
                           RAM_9_9_port, IN4 => n3361, IN5 => n2863, QN => 
                           n2290);
   U2428 : AOI221X1 port map( IN1 => RAM_8_29_port, IN2 => n3417, IN3 => 
                           RAM_9_29_port, IN4 => n3362, IN5 => n2943, QN => 
                           n2282);
   U2429 : AOI221X1 port map( IN1 => RAM_8_63_port, IN2 => n3416, IN3 => 
                           RAM_9_63_port, IN4 => n3368, IN5 => n3079, QN => 
                           n2475);
   U2430 : AOI221X1 port map( IN1 => RAM_8_70_port, IN2 => n3426, IN3 => 
                           RAM_9_70_port, IN4 => n3360, IN5 => n3107, QN => 
                           n2278);
   U2431 : AOI221X1 port map( IN1 => RAM_8_49_port, IN2 => n3423, IN3 => 
                           RAM_9_49_port, IN4 => n3366, IN5 => n3023, QN => 
                           n2606);
   U2432 : AOI221X1 port map( IN1 => RAM_8_116_port, IN2 => n3426, IN3 => 
                           RAM_9_116_port, IN4 => n3364, IN5 => n3295, QN => 
                           n2393);
   U2433 : AOI221X1 port map( IN1 => RAM_8_54_port, IN2 => n3422, IN3 => 
                           RAM_9_54_port, IN4 => n3370, IN5 => n3043, QN => 
                           n2382);
   U2434 : AOI221X1 port map( IN1 => RAM_8_77_port, IN2 => n3422, IN3 => 
                           RAM_9_77_port, IN4 => n3368, IN5 => n3135, QN => 
                           n2294);
   U2435 : AOI221X1 port map( IN1 => RAM_8_64_port, IN2 => n3425, IN3 => 
                           RAM_9_64_port, IN4 => n3367, IN5 => n3083, QN => 
                           n2378);
   U2436 : AOI221X1 port map( IN1 => RAM_8_62_port, IN2 => n3418, IN3 => 
                           RAM_9_62_port, IN4 => n3370, IN5 => n3075, QN => 
                           n2219);
   U2437 : AOI221X1 port map( IN1 => RAM_8_5_port, IN2 => n3419, IN3 => 
                           RAM_9_5_port, IN4 => n3365, IN5 => n2847, QN => 
                           n2802);
   U2438 : AOI221X1 port map( IN1 => RAM_8_76_port, IN2 => n3416, IN3 => 
                           RAM_9_76_port, IN4 => n3366, IN5 => n3131, QN => 
                           n2714);
   U2439 : AOI221X1 port map( IN1 => RAM_8_107_port, IN2 => n3422, IN3 => 
                           RAM_9_107_port, IN4 => n3368, IN5 => n3255, QN => 
                           n2710);
   U2440 : AOI221X1 port map( IN1 => RAM_8_50_port, IN2 => n3415, IN3 => 
                           RAM_9_50_port, IN4 => n3361, IN5 => n3027, QN => 
                           n2412);
   U2441 : AOI221X1 port map( IN1 => RAM_8_72_port, IN2 => n3424, IN3 => 
                           RAM_9_72_port, IN4 => n3365, IN5 => n3115, QN => 
                           n2400);
   U2442 : AOI221X1 port map( IN1 => RAM_8_47_port, IN2 => n3424, IN3 => 
                           RAM_9_47_port, IN4 => n3364, IN5 => n3015, QN => 
                           n2462);
   U2443 : AOI221X1 port map( IN1 => RAM_0_122_port, IN2 => n2165, IN3 => 
                           RAM_1_122_port, IN4 => n3390, IN5 => n3321, QN => 
                           n2483);
   U2444 : INVX0 port map( INP => n3348, ZN => n2621);
   U2445 : INVX0 port map( INP => n3348, ZN => n2622);
   U2446 : AO22X2 port map( IN1 => RAM_11_37_port, IN2 => n3451, IN3 => n2650, 
                           IN4 => RAM_10_37_port, Q => n2975);
   U2447 : NOR2X0 port map( IN1 => n3358, IN2 => RAMADDR1(3), QN => n2202);
   U2448 : AND2X2 port map( IN1 => n2709, IN2 => n2505, Q => n3351);
   U2449 : NAND4X0 port map( IN1 => n2203, IN2 => n2204, IN3 => n2205, IN4 => 
                           n2206, QN => RAMDOUT1(41));
   U2450 : AOI221X1 port map( IN1 => RAM_8_41_port, IN2 => n3418, IN3 => 
                           RAM_9_41_port, IN4 => n3367, IN5 => n2991, QN => 
                           n2203);
   U2451 : AOI221X2 port map( IN1 => RAM_12_41_port, IN2 => n2458, IN3 => 
                           RAM_13_41_port, IN4 => n3371, IN5 => n2992, QN => 
                           n2204);
   U2452 : AOI221X1 port map( IN1 => RAM_0_41_port, IN2 => n2169, IN3 => 
                           RAM_1_41_port, IN4 => n3384, IN5 => n2993, QN => 
                           n2205);
   U2453 : AOI221X1 port map( IN1 => RAM_4_41_port, IN2 => n3407, IN3 => 
                           RAM_5_41_port, IN4 => n3400, IN5 => n2994, QN => 
                           n2206);
   U2454 : NAND4X0 port map( IN1 => n2207, IN2 => n2208, IN3 => n2209, IN4 => 
                           n2210, QN => RAMDOUT1(44));
   U2455 : AOI221X1 port map( IN1 => RAM_12_44_port, IN2 => n2456, IN3 => n3380
                           , IN4 => RAM_13_44_port, IN5 => n3004, QN => n2208);
   U2456 : AOI221X1 port map( IN1 => RAM_0_44_port, IN2 => n2160, IN3 => 
                           RAM_1_44_port, IN4 => n2492, IN5 => n3005, QN => 
                           n2209);
   U2457 : AOI221X2 port map( IN1 => RAM_4_44_port, IN2 => n3408, IN3 => 
                           RAM_5_44_port, IN4 => n3398, IN5 => n3006, QN => 
                           n2210);
   U2458 : AOI221X1 port map( IN1 => RAM_8_34_port, IN2 => n3419, IN3 => 
                           RAM_9_34_port, IN4 => n3364, IN5 => n2963, QN => 
                           n2566);
   U2459 : AOI221X1 port map( IN1 => RAM_0_117_port, IN2 => n2167, IN3 => 
                           RAM_1_117_port, IN4 => n3384, IN5 => n3301, QN => 
                           n2264);
   U2460 : AOI221X1 port map( IN1 => RAM_0_87_port, IN2 => n2165, IN3 => 
                           RAM_1_87_port, IN4 => n2121, IN5 => n3177, QN => 
                           n2434);
   U2461 : AOI221X1 port map( IN1 => RAM_0_96_port, IN2 => n2159, IN3 => 
                           RAM_1_96_port, IN4 => n3385, IN5 => n3213, QN => 
                           n2276);
   U2462 : AOI221X1 port map( IN1 => RAM_0_75_port, IN2 => n2172, IN3 => 
                           RAM_1_75_port, IN4 => n3383, IN5 => n3129, QN => 
                           n2246);
   U2463 : AOI221X1 port map( IN1 => RAM_0_62_port, IN2 => n2162, IN3 => 
                           RAM_1_62_port, IN4 => n3382, IN5 => n3077, QN => 
                           n2221);
   U2464 : AOI221X1 port map( IN1 => RAM_0_39_port, IN2 => n2169, IN3 => 
                           RAM_1_39_port, IN4 => n2157, IN5 => n2985, QN => 
                           n2572);
   U2465 : AOI221X1 port map( IN1 => RAM_0_31_port, IN2 => n2163, IN3 => 
                           RAM_1_31_port, IN4 => n3388, IN5 => n2953, QN => 
                           n2304);
   U2466 : AOI221X1 port map( IN1 => RAM_0_70_port, IN2 => n2166, IN3 => 
                           RAM_1_70_port, IN4 => n3388, IN5 => n3109, QN => 
                           n2280);
   U2467 : AOI221X1 port map( IN1 => RAM_0_119_port, IN2 => n2158, IN3 => 
                           RAM_1_119_port, IN4 => n2157, IN5 => n3309, QN => 
                           n2240);
   U2468 : AOI221X1 port map( IN1 => RAM_0_42_port, IN2 => n2169, IN3 => 
                           RAM_1_42_port, IN4 => n2492, IN5 => n2997, QN => 
                           n2564);
   U2469 : NAND4X0 port map( IN1 => n2211, IN2 => n2212, IN3 => n2213, IN4 => 
                           n2214, QN => RAMDOUT1(43));
   U2470 : AOI221X1 port map( IN1 => RAM_8_43_port, IN2 => n3424, IN3 => 
                           RAM_9_43_port, IN4 => n3360, IN5 => n2999, QN => 
                           n2211);
   U2471 : AOI221X2 port map( IN1 => RAM_12_43_port, IN2 => n2456, IN3 => 
                           RAM_13_43_port, IN4 => n3375, IN5 => n3000, QN => 
                           n2212);
   U2472 : AOI221X1 port map( IN1 => RAM_0_43_port, IN2 => n2171, IN3 => 
                           RAM_1_43_port, IN4 => n3388, IN5 => n3001, QN => 
                           n2213);
   U2473 : AOI221X1 port map( IN1 => RAM_4_43_port, IN2 => n3407, IN3 => 
                           RAM_5_43_port, IN4 => n3395, IN5 => n3002, QN => 
                           n2214);
   U2474 : AOI221X1 port map( IN1 => RAM_0_86_port, IN2 => n2159, IN3 => 
                           RAM_1_86_port, IN4 => n2492, IN5 => n3173, QN => 
                           n2272);
   U2475 : AOI221X1 port map( IN1 => RAM_0_29_port, IN2 => n2169, IN3 => 
                           RAM_1_29_port, IN4 => n3390, IN5 => n2945, QN => 
                           n2284);
   U2476 : NAND4X0 port map( IN1 => n2215, IN2 => n2216, IN3 => n2217, IN4 => 
                           n2218, QN => RAMDOUT1(99));
   U2477 : AOI221X2 port map( IN1 => RAM_8_99_port, IN2 => n3418, IN3 => 
                           RAM_9_99_port, IN4 => n3369, IN5 => n3223, QN => 
                           n2215);
   U2478 : AOI221X2 port map( IN1 => RAM_4_99_port, IN2 => n3410, IN3 => 
                           RAM_5_99_port, IN4 => n3397, IN5 => n3226, QN => 
                           n2216);
   U2479 : AOI221X2 port map( IN1 => RAM_12_99_port, IN2 => n2453, IN3 => 
                           RAM_13_99_port, IN4 => n3378, IN5 => n3224, QN => 
                           n2218);
   U2480 : AOI221X1 port map( IN1 => RAM_0_72_port, IN2 => n2166, IN3 => 
                           RAM_1_72_port, IN4 => n2157, IN5 => n3117, QN => 
                           n2402);
   U2481 : AOI221X1 port map( IN1 => RAM_4_107_port, IN2 => n3405, IN3 => 
                           RAM_5_107_port, IN4 => n3400, IN5 => n3258, QN => 
                           n2713);
   U2482 : NAND4X0 port map( IN1 => n2219, IN2 => n2220, IN3 => n2221, IN4 => 
                           n2222, QN => RAMDOUT1(62));
   U2483 : AOI221X1 port map( IN1 => RAM_12_62_port, IN2 => n2446, IN3 => n3380
                           , IN4 => RAM_13_62_port, IN5 => n3076, QN => n2220);
   U2484 : AOI221X2 port map( IN1 => RAM_4_62_port, IN2 => n3402, IN3 => 
                           RAM_5_62_port, IN4 => n3401, IN5 => n3078, QN => 
                           n2222);
   U2485 : NAND4X0 port map( IN1 => n2223, IN2 => n2224, IN3 => n2225, IN4 => 
                           n2226, QN => RAMDOUT1(11));
   U2486 : AOI221X1 port map( IN1 => RAM_12_11_port, IN2 => n2453, IN3 => n3374
                           , IN4 => RAM_13_11_port, IN5 => n2872, QN => n2224);
   U2487 : AOI221X1 port map( IN1 => RAM_0_11_port, IN2 => n2167, IN3 => 
                           RAM_1_11_port, IN4 => n3383, IN5 => n2873, QN => 
                           n2225);
   U2488 : AOI221X2 port map( IN1 => RAM_4_11_port, IN2 => n3409, IN3 => 
                           RAM_5_11_port, IN4 => n2495, IN5 => n2874, QN => 
                           n2226);
   U2489 : NAND4X0 port map( IN1 => n2227, IN2 => n2228, IN3 => n2229, IN4 => 
                           n2230, QN => RAMDOUT1(19));
   U2490 : AOI221X2 port map( IN1 => RAM_8_19_port, IN2 => n3417, IN3 => 
                           RAM_9_19_port, IN4 => n3368, IN5 => n2903, QN => 
                           n2227);
   U2491 : AOI221X1 port map( IN1 => RAM_12_19_port, IN2 => n2452, IN3 => n3375
                           , IN4 => RAM_13_19_port, IN5 => n2904, QN => n2228);
   U2492 : AOI221X1 port map( IN1 => RAM_0_19_port, IN2 => n2164, IN3 => 
                           RAM_1_19_port, IN4 => n3384, IN5 => n2905, QN => 
                           n2229);
   U2493 : AOI221X2 port map( IN1 => RAM_4_19_port, IN2 => n3403, IN3 => 
                           RAM_5_19_port, IN4 => n2494, IN5 => n2906, QN => 
                           n2230);
   U2494 : INVX0 port map( INP => n2499, ZN => n2231);
   U2495 : NAND4X0 port map( IN1 => n2232, IN2 => n2233, IN3 => n2234, IN4 => 
                           n2235, QN => RAMDOUT1(55));
   U2496 : AOI221X1 port map( IN1 => RAM_12_55_port, IN2 => n2448, IN3 => n3373
                           , IN4 => RAM_13_55_port, IN5 => n3048, QN => n2233);
   U2497 : AOI221X2 port map( IN1 => RAM_4_55_port, IN2 => n3409, IN3 => 
                           RAM_5_55_port, IN4 => n3398, IN5 => n3050, QN => 
                           n2235);
   U2498 : NAND4X0 port map( IN1 => n2236, IN2 => n2238, IN3 => n2237, IN4 => 
                           n2239, QN => RAMDOUT1(85));
   U2499 : AOI221X2 port map( IN1 => RAM_12_85_port, IN2 => n2454, IN3 => 
                           RAM_13_85_port, IN4 => n3376, IN5 => n3168, QN => 
                           n2237);
   U2500 : AOI221X2 port map( IN1 => RAM_4_85_port, IN2 => n3409, IN3 => 
                           RAM_5_85_port, IN4 => n2494, IN5 => n3170, QN => 
                           n2239);
   U2501 : NAND4X0 port map( IN1 => n2240, IN2 => n2241, IN3 => n2242, IN4 => 
                           n2243, QN => RAMDOUT1(119));
   U2502 : AOI221X2 port map( IN1 => RAM_12_119_port, IN2 => n2447, IN3 => 
                           RAM_13_119_port, IN4 => n3372, IN5 => n3308, QN => 
                           n2241);
   U2503 : NAND4X0 port map( IN1 => n2246, IN2 => n2244, IN3 => n2245, IN4 => 
                           n2247, QN => RAMDOUT1(75));
   U2504 : AOI221X2 port map( IN1 => RAM_12_75_port, IN2 => n2453, IN3 => 
                           RAM_13_75_port, IN4 => n3378, IN5 => n3128, QN => 
                           n2245);
   U2505 : AOI221X2 port map( IN1 => RAM_4_75_port, IN2 => n3409, IN3 => 
                           RAM_5_75_port, IN4 => n3392, IN5 => n3130, QN => 
                           n2247);
   U2506 : NBUFFX2 port map( INP => RAMDIN1(22), Z => n2248);
   U2507 : NBUFFX2 port map( INP => RAMDIN1(22), Z => n2249);
   U2508 : NAND4X0 port map( IN1 => n2252, IN2 => n2251, IN3 => n2250, IN4 => 
                           n2253, QN => RAMDOUT1(89));
   U2509 : AOI221X1 port map( IN1 => RAM_8_89_port, IN2 => n3423, IN3 => 
                           RAM_9_89_port, IN4 => n3365, IN5 => n3183, QN => 
                           n2250);
   U2510 : AOI221X2 port map( IN1 => RAM_4_89_port, IN2 => n3406, IN3 => 
                           RAM_5_89_port, IN4 => n3395, IN5 => n3186, QN => 
                           n2253);
   U2511 : NAND4X0 port map( IN1 => n2254, IN2 => n2255, IN3 => n2256, IN4 => 
                           n2257, QN => RAMDOUT1(83));
   U2512 : AOI221X1 port map( IN1 => RAM_8_83_port, IN2 => n3425, IN3 => 
                           RAM_9_83_port, IN4 => n3367, IN5 => n3159, QN => 
                           n2254);
   U2513 : AOI221X2 port map( IN1 => RAM_4_83_port, IN2 => n3403, IN3 => 
                           RAM_5_83_port, IN4 => n3401, IN5 => n3162, QN => 
                           n2257);
   U2514 : NAND4X0 port map( IN1 => n2258, IN2 => n2260, IN3 => n2259, IN4 => 
                           n2261, QN => RAMDOUT1(111));
   U2515 : AOI221X1 port map( IN1 => RAM_8_111_port, IN2 => n3422, IN3 => 
                           RAM_9_111_port, IN4 => n3370, IN5 => n3271, QN => 
                           n2258);
   U2516 : AOI221X2 port map( IN1 => RAM_12_111_port, IN2 => n2447, IN3 => 
                           RAM_13_111_port, IN4 => n3373, IN5 => n3272, QN => 
                           n2259);
   U2517 : AOI221X1 port map( IN1 => RAM_0_111_port, IN2 => n2165, IN3 => 
                           RAM_1_111_port, IN4 => n3384, IN5 => n3273, QN => 
                           n2260);
   U2518 : NAND4X0 port map( IN1 => n2262, IN2 => n2263, IN3 => n2264, IN4 => 
                           n2265, QN => RAMDOUT1(117));
   U2519 : AOI221X2 port map( IN1 => RAM_12_117_port, IN2 => n2446, IN3 => 
                           RAM_13_117_port, IN4 => n3373, IN5 => n3300, QN => 
                           n2263);
   U2520 : AOI221X2 port map( IN1 => RAM_4_117_port, IN2 => n3402, IN3 => 
                           RAM_5_117_port, IN4 => n3399, IN5 => n3302, QN => 
                           n2265);
   U2521 : NAND4X0 port map( IN1 => n2266, IN2 => n2267, IN3 => n2268, IN4 => 
                           n2269, QN => RAMDOUT1(90));
   U2522 : AOI221X2 port map( IN1 => RAM_12_90_port, IN2 => n2452, IN3 => 
                           RAM_13_90_port, IN4 => n3371, IN5 => n3188, QN => 
                           n2267);
   U2523 : AOI221X1 port map( IN1 => RAM_0_90_port, IN2 => n2168, IN3 => 
                           RAM_1_90_port, IN4 => n3390, IN5 => n3189, QN => 
                           n2268);
   U2524 : AOI221X2 port map( IN1 => RAM_4_90_port, IN2 => n3402, IN3 => 
                           RAM_5_90_port, IN4 => n3397, IN5 => n3190, QN => 
                           n2269);
   U2525 : NAND4X0 port map( IN1 => n2270, IN2 => n2271, IN3 => n2272, IN4 => 
                           n2273, QN => RAMDOUT1(86));
   U2526 : AOI221X1 port map( IN1 => RAM_8_86_port, IN2 => n3418, IN3 => 
                           RAM_9_86_port, IN4 => n3361, IN5 => n3171, QN => 
                           n2270);
   U2527 : AOI221X2 port map( IN1 => RAM_12_86_port, IN2 => n2445, IN3 => 
                           RAM_13_86_port, IN4 => n3375, IN5 => n3172, QN => 
                           n2271);
   U2528 : AOI221X2 port map( IN1 => RAM_4_86_port, IN2 => n3405, IN3 => 
                           RAM_5_86_port, IN4 => n3398, IN5 => n3174, QN => 
                           n2273);
   U2529 : NAND4X0 port map( IN1 => n2274, IN2 => n2275, IN3 => n2276, IN4 => 
                           n2277, QN => RAMDOUT1(96));
   U2530 : AOI221X2 port map( IN1 => RAM_12_96_port, IN2 => n2448, IN3 => 
                           RAM_13_96_port, IN4 => n3373, IN5 => n3212, QN => 
                           n2275);
   U2531 : AOI221X2 port map( IN1 => RAM_4_96_port, IN2 => n3408, IN3 => 
                           RAM_5_96_port, IN4 => n3397, IN5 => n3214, QN => 
                           n2277);
   U2532 : NAND4X0 port map( IN1 => n2280, IN2 => n2279, IN3 => n2278, IN4 => 
                           n2281, QN => RAMDOUT1(70));
   U2533 : AOI221X2 port map( IN1 => RAM_12_70_port, IN2 => n2447, IN3 => 
                           RAM_13_70_port, IN4 => n2490, IN5 => n3108, QN => 
                           n2279);
   U2534 : AOI221X2 port map( IN1 => RAM_4_70_port, IN2 => n3406, IN3 => 
                           RAM_5_70_port, IN4 => n2495, IN5 => n3110, QN => 
                           n2281);
   U2535 : NAND4X0 port map( IN1 => n2282, IN2 => n2283, IN3 => n2284, IN4 => 
                           n2285, QN => RAMDOUT1(29));
   U2536 : AOI221X2 port map( IN1 => RAM_12_29_port, IN2 => n2449, IN3 => 
                           RAM_13_29_port, IN4 => n2489, IN5 => n2944, QN => 
                           n2283);
   U2537 : AOI221X2 port map( IN1 => RAM_4_29_port, IN2 => n3406, IN3 => 
                           RAM_5_29_port, IN4 => n3398, IN5 => n2946, QN => 
                           n2285);
   U2538 : NAND4X0 port map( IN1 => n2286, IN2 => n2287, IN3 => n2288, IN4 => 
                           n2289, QN => RAMDOUT1(60));
   U2539 : AOI221X2 port map( IN1 => RAM_12_60_port, IN2 => n2458, IN3 => 
                           RAM_13_60_port, IN4 => n3376, IN5 => n3068, QN => 
                           n2287);
   U2540 : AOI221X2 port map( IN1 => RAM_0_60_port, IN2 => n2164, IN3 => 
                           RAM_1_60_port, IN4 => n2492, IN5 => n3069, QN => 
                           n2288);
   U2541 : AOI221X2 port map( IN1 => RAM_4_60_port, IN2 => n3404, IN3 => 
                           RAM_5_60_port, IN4 => n3399, IN5 => n3070, QN => 
                           n2289);
   U2542 : NAND4X0 port map( IN1 => n2290, IN2 => n2291, IN3 => n2292, IN4 => 
                           n2293, QN => RAMDOUT1(9));
   U2543 : AOI221X2 port map( IN1 => RAM_12_9_port, IN2 => n2456, IN3 => 
                           RAM_13_9_port, IN4 => n3377, IN5 => n2864, QN => 
                           n2291);
   U2544 : AOI221X2 port map( IN1 => RAM_4_9_port, IN2 => n3406, IN3 => 
                           RAM_5_9_port, IN4 => n3391, IN5 => n2866, QN => 
                           n2293);
   U2545 : NAND4X0 port map( IN1 => n2294, IN2 => n2295, IN3 => n2296, IN4 => 
                           n2297, QN => RAMDOUT1(77));
   U2546 : AOI221X2 port map( IN1 => RAM_12_77_port, IN2 => n2452, IN3 => 
                           RAM_13_77_port, IN4 => n3380, IN5 => n3136, QN => 
                           n2295);
   U2547 : AOI221X2 port map( IN1 => RAM_4_77_port, IN2 => n3448, IN3 => 
                           RAM_5_77_port, IN4 => n3391, IN5 => n3138, QN => 
                           n2297);
   U2548 : NAND4X0 port map( IN1 => n2298, IN2 => n2299, IN3 => n2300, IN4 => 
                           n2301, QN => RAMDOUT1(10));
   U2549 : AOI221X2 port map( IN1 => RAM_12_10_port, IN2 => n2459, IN3 => 
                           RAM_13_10_port, IN4 => n3378, IN5 => n2868, QN => 
                           n2299);
   U2550 : AOI221X2 port map( IN1 => RAM_4_10_port, IN2 => n3407, IN3 => 
                           RAM_5_10_port, IN4 => n3394, IN5 => n2870, QN => 
                           n2301);
   U2551 : NAND4X0 port map( IN1 => n2302, IN2 => n2303, IN3 => n2304, IN4 => 
                           n2305, QN => RAMDOUT1(31));
   U2552 : AOI221X2 port map( IN1 => RAM_8_31_port, IN2 => n3425, IN3 => 
                           RAM_9_31_port, IN4 => n3360, IN5 => n2951, QN => 
                           n2302);
   U2553 : AOI221X2 port map( IN1 => RAM_12_31_port, IN2 => n2451, IN3 => 
                           RAM_13_31_port, IN4 => n3376, IN5 => n2952, QN => 
                           n2303);
   U2554 : AOI221X2 port map( IN1 => RAM_4_31_port, IN2 => n3410, IN3 => 
                           RAM_5_31_port, IN4 => n2495, IN5 => n2954, QN => 
                           n2305);
   U2555 : NAND4X0 port map( IN1 => n2306, IN2 => n2307, IN3 => n2308, IN4 => 
                           n2309, QN => RAMDOUT1(97));
   U2556 : AOI221X2 port map( IN1 => RAM_12_97_port, IN2 => n2454, IN3 => 
                           RAM_13_97_port, IN4 => n3381, IN5 => n3216, QN => 
                           n2307);
   U2557 : AOI221X2 port map( IN1 => RAM_4_97_port, IN2 => n3406, IN3 => 
                           RAM_5_97_port, IN4 => n3396, IN5 => n3218, QN => 
                           n2309);
   U2558 : NAND4X0 port map( IN1 => n2310, IN2 => n2311, IN3 => n2312, IN4 => 
                           n2313, QN => RAMDOUT1(103));
   U2559 : AOI221X1 port map( IN1 => RAM_8_103_port, IN2 => n3421, IN3 => 
                           RAM_9_103_port, IN4 => n3370, IN5 => n3239, QN => 
                           n2310);
   U2560 : AOI221X2 port map( IN1 => RAM_12_103_port, IN2 => n2449, IN3 => 
                           RAM_13_103_port, IN4 => n3377, IN5 => n3240, QN => 
                           n2311);
   U2561 : AOI221X1 port map( IN1 => RAM_0_103_port, IN2 => n2167, IN3 => 
                           RAM_1_103_port, IN4 => n2157, IN5 => n3241, QN => 
                           n2312);
   U2562 : AOI221X2 port map( IN1 => RAM_4_103_port, IN2 => n3448, IN3 => 
                           RAM_5_103_port, IN4 => n3396, IN5 => n3242, QN => 
                           n2313);
   U2563 : NAND4X0 port map( IN1 => n2314, IN2 => n2315, IN3 => n2316, IN4 => 
                           n2317, QN => RAMDOUT1(7));
   U2564 : AOI221X2 port map( IN1 => RAM_12_7_port, IN2 => n2455, IN3 => 
                           RAM_13_7_port, IN4 => n3379, IN5 => n2856, QN => 
                           n2315);
   U2565 : AOI221X2 port map( IN1 => RAM_4_7_port, IN2 => n3404, IN3 => 
                           RAM_5_7_port, IN4 => n3394, IN5 => n2858, QN => 
                           n2317);
   U2566 : AO22X2 port map( IN1 => RAM_11_45_port, IN2 => n2501, IN3 => n2662, 
                           IN4 => RAM_10_45_port, Q => n3007);
   U2567 : AO22X2 port map( IN1 => RAM_11_79_port, IN2 => n2498, IN3 => n2112, 
                           IN4 => RAM_10_79_port, Q => n3143);
   U2568 : AO22X2 port map( IN1 => RAM_11_66_port, IN2 => n3450, IN3 => n2650, 
                           IN4 => RAM_10_66_port, Q => n3091);
   U2569 : AO22X2 port map( IN1 => RAM_11_63_port, IN2 => n2466, IN3 => 
                           RAM_10_63_port, IN4 => n2666, Q => n3079);
   U2570 : AO22X2 port map( IN1 => RAM_11_42_port, IN2 => n3452, IN3 => 
                           RAM_10_42_port, IN4 => n2664, Q => n2995);
   U2571 : AO22X2 port map( IN1 => RAM_11_47_port, IN2 => n3461, IN3 => n2112, 
                           IN4 => RAM_10_47_port, Q => n3015);
   U2572 : AO22X2 port map( IN1 => RAM_11_32_port, IN2 => n3462, IN3 => 
                           RAM_10_32_port, IN4 => n2661, Q => n2955);
   U2573 : AO22X2 port map( IN1 => RAM_11_67_port, IN2 => n2498, IN3 => 
                           RAM_10_67_port, IN4 => n2661, Q => n3095);
   U2574 : AO22X2 port map( IN1 => RAM_11_56_port, IN2 => n3451, IN3 => n2461, 
                           IN4 => RAM_10_56_port, Q => n3051);
   U2575 : AND2X4 port map( IN1 => n2797, IN2 => n2821, Q => n2318);
   U2576 : AND2X4 port map( IN1 => n2797, IN2 => n2821, Q => n2319);
   U2577 : NBUFFX2 port map( INP => n2318, Z => n2320);
   U2578 : DELLN1X2 port map( INP => n2318, Z => n2321);
   U2579 : NBUFFX2 port map( INP => n2318, Z => n2322);
   U2580 : DELLN1X2 port map( INP => n2318, Z => n2323);
   U2581 : NBUFFX2 port map( INP => n2319, Z => n2325);
   U2582 : NBUFFX2 port map( INP => n2319, Z => n2326);
   U2583 : NBUFFX2 port map( INP => n2319, Z => n2327);
   U2584 : NBUFFX2 port map( INP => n2319, Z => n2328);
   U2585 : NBUFFX2 port map( INP => n2319, Z => n2329);
   U2586 : NBUFFX2 port map( INP => n3343, Z => n2330);
   U2587 : NBUFFX2 port map( INP => n3343, Z => n2331);
   U2588 : NBUFFX2 port map( INP => n3343, Z => n2332);
   U2589 : NBUFFX2 port map( INP => n3343, Z => n2333);
   U2590 : NBUFFX2 port map( INP => n3343, Z => n2334);
   U2591 : NBUFFX2 port map( INP => n2748, Z => n2335);
   U2592 : NBUFFX2 port map( INP => n2748, Z => n2336);
   U2593 : NBUFFX2 port map( INP => n2748, Z => n2337);
   U2594 : NBUFFX2 port map( INP => n2748, Z => n2338);
   U2595 : NBUFFX2 port map( INP => n2748, Z => n2339);
   U2596 : INVX0 port map( INP => n2509, ZN => n2340);
   U2597 : AND2X1 port map( IN1 => n5615, IN2 => RAMADDR1(1), Q => n2828);
   U2598 : NAND4X0 port map( IN1 => n2341, IN2 => n2342, IN3 => n2343, IN4 => 
                           n2344, QN => RAMDOUT1(127));
   U2599 : AOI221X2 port map( IN1 => RAM_12_127_port, IN2 => n2452, IN3 => 
                           RAM_13_127_port, IN4 => n3377, IN5 => n3345, QN => 
                           n2342);
   U2600 : AOI221X2 port map( IN1 => RAM_0_127_port, IN2 => n2168, IN3 => 
                           RAM_1_127_port, IN4 => n3383, IN5 => n3350, QN => 
                           n2343);
   U2601 : NAND4X0 port map( IN1 => n2345, IN2 => n2346, IN3 => n2347, IN4 => 
                           n2348, QN => RAMDOUT1(40));
   U2602 : AOI221X2 port map( IN1 => RAM_12_40_port, IN2 => n2450, IN3 => 
                           RAM_13_40_port, IN4 => n3374, IN5 => n2988, QN => 
                           n2346);
   U2603 : AOI221X1 port map( IN1 => RAM_0_40_port, IN2 => n2170, IN3 => 
                           RAM_1_40_port, IN4 => n3387, IN5 => n2989, QN => 
                           n2347);
   U2604 : AOI221X2 port map( IN1 => RAM_4_40_port, IN2 => n3410, IN3 => 
                           RAM_5_40_port, IN4 => n3394, IN5 => n2990, QN => 
                           n2348);
   U2605 : NAND4X0 port map( IN1 => n2349, IN2 => n2350, IN3 => n2351, IN4 => 
                           n2352, QN => RAMDOUT1(36));
   U2606 : AOI221X2 port map( IN1 => RAM_12_36_port, IN2 => n2455, IN3 => 
                           RAM_13_36_port, IN4 => n3377, IN5 => n2972, QN => 
                           n2350);
   U2607 : AOI221X1 port map( IN1 => RAM_0_36_port, IN2 => n2164, IN3 => 
                           RAM_1_36_port, IN4 => n2492, IN5 => n2973, QN => 
                           n2351);
   U2608 : AOI221X2 port map( IN1 => RAM_4_36_port, IN2 => n3407, IN3 => 
                           RAM_5_36_port, IN4 => n3393, IN5 => n2974, QN => 
                           n2352);
   U2609 : NAND4X0 port map( IN1 => n2353, IN2 => n2354, IN3 => n2355, IN4 => 
                           n2356, QN => RAMDOUT1(1));
   U2610 : AOI221X2 port map( IN1 => RAM_12_1_port, IN2 => n2458, IN3 => 
                           RAM_13_1_port, IN4 => n2489, IN5 => n2832, QN => 
                           n2354);
   U2611 : AOI221X1 port map( IN1 => RAM_0_1_port, IN2 => n2163, IN3 => 
                           RAM_1_1_port, IN4 => n3387, IN5 => n2833, QN => 
                           n2355);
   U2612 : AOI221X2 port map( IN1 => RAM_4_1_port, IN2 => n3402, IN3 => 
                           RAM_5_1_port, IN4 => n3398, IN5 => n2834, QN => 
                           n2356);
   U2613 : NAND4X0 port map( IN1 => n2357, IN2 => n2358, IN3 => n2359, IN4 => 
                           n2360, QN => RAMDOUT1(35));
   U2614 : AOI221X2 port map( IN1 => RAM_12_35_port, IN2 => n2445, IN3 => 
                           RAM_13_35_port, IN4 => n2490, IN5 => n2968, QN => 
                           n2358);
   U2615 : NAND4X0 port map( IN1 => n2361, IN2 => n2362, IN3 => n2363, IN4 => 
                           n2364, QN => RAMDOUT1(58));
   U2616 : AOI221X2 port map( IN1 => RAM_12_58_port, IN2 => n2454, IN3 => 
                           RAM_13_58_port, IN4 => n3371, IN5 => n3060, QN => 
                           n2362);
   U2617 : AOI221X2 port map( IN1 => RAM_4_58_port, IN2 => n3409, IN3 => 
                           RAM_5_58_port, IN4 => n2494, IN5 => n3062, QN => 
                           n2364);
   U2618 : NAND4X0 port map( IN1 => n2365, IN2 => n2366, IN3 => n2367, IN4 => 
                           n2368, QN => RAMDOUT1(12));
   U2619 : AOI221X2 port map( IN1 => RAM_12_12_port, IN2 => n2451, IN3 => 
                           RAM_13_12_port, IN4 => n3379, IN5 => n2876, QN => 
                           n2366);
   U2620 : AOI221X1 port map( IN1 => RAM_0_12_port, IN2 => n2168, IN3 => 
                           RAM_1_12_port, IN4 => n3386, IN5 => n2877, QN => 
                           n2367);
   U2621 : AOI221X2 port map( IN1 => RAM_4_12_port, IN2 => n3403, IN3 => 
                           RAM_5_12_port, IN4 => n2494, IN5 => n2878, QN => 
                           n2368);
   U2622 : NAND4X0 port map( IN1 => n2369, IN2 => n2370, IN3 => n2371, IN4 => 
                           n2372, QN => RAMDOUT1(105));
   U2623 : AOI221X2 port map( IN1 => RAM_12_105_port, IN2 => n2451, IN3 => 
                           RAM_13_105_port, IN4 => n3375, IN5 => n3248, QN => 
                           n2370);
   U2624 : AOI221X2 port map( IN1 => RAM_4_105_port, IN2 => n3404, IN3 => 
                           RAM_5_105_port, IN4 => n3392, IN5 => n3250, QN => 
                           n2372);
   U2625 : INVX0 port map( INP => n2647, ZN => n2373);
   U2626 : NAND4X0 port map( IN1 => n2374, IN2 => n2375, IN3 => n2376, IN4 => 
                           n2377, QN => RAMDOUT1(73));
   U2627 : AOI221X2 port map( IN1 => RAM_12_73_port, IN2 => n2457, IN3 => 
                           RAM_13_73_port, IN4 => n3381, IN5 => n3120, QN => 
                           n2375);
   U2628 : AOI221X2 port map( IN1 => RAM_4_73_port, IN2 => n3402, IN3 => 
                           RAM_5_73_port, IN4 => n3396, IN5 => n3122, QN => 
                           n2377);
   U2629 : NAND4X0 port map( IN1 => n2378, IN2 => n2379, IN3 => n2380, IN4 => 
                           n2381, QN => RAMDOUT1(64));
   U2630 : AOI221X1 port map( IN1 => RAM_12_64_port, IN2 => n2446, IN3 => 
                           RAM_13_64_port, IN4 => n3378, IN5 => n3084, QN => 
                           n2379);
   U2631 : AOI221X1 port map( IN1 => RAM_0_64_port, IN2 => n2161, IN3 => 
                           RAM_1_64_port, IN4 => n3382, IN5 => n3085, QN => 
                           n2380);
   U2632 : AOI221X2 port map( IN1 => RAM_4_64_port, IN2 => n3448, IN3 => 
                           RAM_5_64_port, IN4 => n3393, IN5 => n3086, QN => 
                           n2381);
   U2633 : NAND4X0 port map( IN1 => n2382, IN2 => n2383, IN3 => n2384, IN4 => 
                           n2385, QN => RAMDOUT1(54));
   U2634 : AOI221X2 port map( IN1 => RAM_12_54_port, IN2 => n2449, IN3 => 
                           RAM_13_54_port, IN4 => n3372, IN5 => n3044, QN => 
                           n2383);
   U2635 : AOI221X1 port map( IN1 => RAM_0_54_port, IN2 => n2164, IN3 => 
                           RAM_1_54_port, IN4 => n2121, IN5 => n3045, QN => 
                           n2384);
   U2636 : AOI221X2 port map( IN1 => RAM_4_54_port, IN2 => n3403, IN3 => 
                           RAM_5_54_port, IN4 => n3392, IN5 => n3046, QN => 
                           n2385);
   U2637 : NAND4X0 port map( IN1 => n2386, IN2 => n2387, IN3 => n2388, IN4 => 
                           n2389, QN => RAMDOUT1(65));
   U2638 : AOI221X2 port map( IN1 => RAM_12_65_port, IN2 => n2448, IN3 => 
                           RAM_13_65_port, IN4 => n3371, IN5 => n3088, QN => 
                           n2387);
   U2639 : AOI221X1 port map( IN1 => RAM_0_65_port, IN2 => n2167, IN3 => 
                           RAM_1_65_port, IN4 => n3388, IN5 => n3089, QN => 
                           n2388);
   U2640 : AOI221X2 port map( IN1 => RAM_4_65_port, IN2 => n3407, IN3 => 
                           RAM_5_65_port, IN4 => n3394, IN5 => n3090, QN => 
                           n2389);
   U2641 : NAND4X0 port map( IN1 => n2390, IN2 => n2391, IN3 => n2392, IN4 => 
                           n2393, QN => RAMDOUT1(116));
   U2642 : AOI221X2 port map( IN1 => RAM_4_116_port, IN2 => n3406, IN3 => 
                           RAM_5_116_port, IN4 => n3393, IN5 => n3298, QN => 
                           n2390);
   U2643 : AOI221X2 port map( IN1 => RAM_12_116_port, IN2 => n2456, IN3 => 
                           RAM_13_116_port, IN4 => n3374, IN5 => n3296, QN => 
                           n2391);
   U2644 : AOI221X2 port map( IN1 => RAM_0_116_port, IN2 => n2169, IN3 => 
                           RAM_1_116_port, IN4 => n3389, IN5 => n3297, QN => 
                           n2392);
   U2645 : AOI221X1 port map( IN1 => RAM_0_49_port, IN2 => n2168, IN3 => 
                           RAM_1_49_port, IN4 => n3383, IN5 => n3025, QN => 
                           n2608);
   U2646 : AOI221X1 port map( IN1 => RAM_0_34_port, IN2 => n2163, IN3 => 
                           RAM_1_34_port, IN4 => n3385, IN5 => n2965, QN => 
                           n2568);
   U2647 : AOI221X1 port map( IN1 => RAM_0_118_port, IN2 => n2172, IN3 => 
                           RAM_1_118_port, IN4 => n3387, IN5 => n3305, QN => 
                           n2600);
   U2648 : AOI221X1 port map( IN1 => RAM_0_78_port, IN2 => n2173, IN3 => 
                           RAM_1_78_port, IN4 => n3388, IN5 => n3141, QN => 
                           n2678);
   U2649 : AOI221X1 port map( IN1 => RAM_0_109_port, IN2 => n2160, IN3 => 
                           RAM_1_109_port, IN4 => n3383, IN5 => n3265, QN => 
                           n2438);
   U2650 : AOI221X1 port map( IN1 => RAM_0_56_port, IN2 => n2163, IN3 => 
                           RAM_1_56_port, IN4 => n3383, IN5 => n3053, QN => 
                           n2604);
   U2651 : AOI221X1 port map( IN1 => RAM_0_15_port, IN2 => n2166, IN3 => 
                           RAM_1_15_port, IN4 => n3384, IN5 => n2889, QN => 
                           n2422);
   U2652 : AOI221X1 port map( IN1 => RAM_0_114_port, IN2 => n2158, IN3 => 
                           RAM_1_114_port, IN4 => n3382, IN5 => n3289, QN => 
                           n2596);
   U2653 : INVX0 port map( INP => n2511, ZN => n2394);
   U2654 : INVX0 port map( INP => n3354, ZN => n2511);
   U2655 : NAND4X0 port map( IN1 => n2395, IN2 => n2396, IN3 => n2397, IN4 => 
                           n2398, QN => RAMDOUT1(91));
   U2656 : AOI221X1 port map( IN1 => RAM_8_91_port, IN2 => n3418, IN3 => 
                           RAM_9_91_port, IN4 => n3370, IN5 => n3191, QN => 
                           n2395);
   U2657 : AOI221X2 port map( IN1 => RAM_12_91_port, IN2 => n2451, IN3 => 
                           RAM_13_91_port, IN4 => n3374, IN5 => n3192, QN => 
                           n2396);
   U2658 : AOI221X1 port map( IN1 => RAM_0_91_port, IN2 => n2168, IN3 => 
                           RAM_1_91_port, IN4 => n3390, IN5 => n3193, QN => 
                           n2397);
   U2659 : AOI221X2 port map( IN1 => RAM_4_91_port, IN2 => n3408, IN3 => 
                           RAM_5_91_port, IN4 => n3392, IN5 => n3194, QN => 
                           n2398);
   U2660 : IBUFFX16 port map( INP => n2534, ZN => n2399);
   U2661 : INVX0 port map( INP => n3349, ZN => n2536);
   U2662 : NAND4X0 port map( IN1 => n2400, IN2 => n2401, IN3 => n2402, IN4 => 
                           n2403, QN => RAMDOUT1(72));
   U2663 : AOI221X2 port map( IN1 => RAM_12_72_port, IN2 => n2445, IN3 => 
                           RAM_13_72_port, IN4 => n3381, IN5 => n3116, QN => 
                           n2401);
   U2664 : AOI221X2 port map( IN1 => RAM_4_72_port, IN2 => n3407, IN3 => 
                           RAM_5_72_port, IN4 => n3396, IN5 => n3118, QN => 
                           n2403);
   U2665 : NAND4X0 port map( IN1 => n2404, IN2 => n2405, IN3 => n2406, IN4 => 
                           n2407, QN => RAMDOUT1(16));
   U2666 : AOI221X2 port map( IN1 => RAM_12_16_port, IN2 => n2460, IN3 => 
                           RAM_13_16_port, IN4 => n3379, IN5 => n2892, QN => 
                           n2405);
   U2667 : AOI221X1 port map( IN1 => RAM_0_16_port, IN2 => n2166, IN3 => 
                           RAM_1_16_port, IN4 => n3386, IN5 => n2893, QN => 
                           n2406);
   U2668 : AOI221X2 port map( IN1 => RAM_4_16_port, IN2 => n3403, IN3 => 
                           RAM_5_16_port, IN4 => n3395, IN5 => n2894, QN => 
                           n2407);
   U2669 : NAND4X0 port map( IN1 => n2408, IN2 => n2409, IN3 => n2410, IN4 => 
                           n2411, QN => RAMDOUT1(18));
   U2670 : AOI221X2 port map( IN1 => RAM_12_18_port, IN2 => n2459, IN3 => 
                           RAM_13_18_port, IN4 => n3372, IN5 => n2900, QN => 
                           n2409);
   U2671 : AOI221X1 port map( IN1 => RAM_0_18_port, IN2 => n2163, IN3 => 
                           RAM_1_18_port, IN4 => n3389, IN5 => n2901, QN => 
                           n2410);
   U2672 : NAND4X0 port map( IN1 => n2412, IN2 => n2413, IN3 => n2414, IN4 => 
                           n2415, QN => RAMDOUT1(50));
   U2673 : AOI221X2 port map( IN1 => RAM_12_50_port, IN2 => n2450, IN3 => 
                           RAM_13_50_port, IN4 => n3381, IN5 => n3028, QN => 
                           n2413);
   U2674 : AOI221X1 port map( IN1 => RAM_0_50_port, IN2 => n2161, IN3 => 
                           RAM_1_50_port, IN4 => n2121, IN5 => n3029, QN => 
                           n2414);
   U2675 : AOI221X2 port map( IN1 => RAM_4_50_port, IN2 => n3407, IN3 => 
                           RAM_5_50_port, IN4 => n3400, IN5 => n3030, QN => 
                           n2415);
   U2676 : NAND4X0 port map( IN1 => n2416, IN2 => n2417, IN3 => n2418, IN4 => 
                           n2419, QN => RAMDOUT1(17));
   U2677 : AOI221X1 port map( IN1 => RAM_12_17_port, IN2 => n2445, IN3 => 
                           RAM_13_17_port, IN4 => n3376, IN5 => n2896, QN => 
                           n2417);
   U2678 : AOI221X1 port map( IN1 => RAM_0_17_port, IN2 => n2167, IN3 => 
                           RAM_1_17_port, IN4 => n3389, IN5 => n2897, QN => 
                           n2418);
   U2679 : AOI221X2 port map( IN1 => RAM_4_17_port, IN2 => n3408, IN3 => 
                           RAM_5_17_port, IN4 => n3396, IN5 => n2898, QN => 
                           n2419);
   U2680 : NAND4X0 port map( IN1 => n2420, IN2 => n2421, IN3 => n2422, IN4 => 
                           n2423, QN => RAMDOUT1(15));
   U2681 : AOI221X2 port map( IN1 => RAM_12_15_port, IN2 => n2453, IN3 => 
                           RAM_13_15_port, IN4 => n3375, IN5 => n2888, QN => 
                           n2421);
   U2682 : AOI221X2 port map( IN1 => RAM_4_15_port, IN2 => n3410, IN3 => 
                           RAM_5_15_port, IN4 => n3401, IN5 => n2890, QN => 
                           n2423);
   U2683 : NAND4X0 port map( IN1 => n2424, IN2 => n2425, IN3 => n2426, IN4 => 
                           n2427, QN => RAMDOUT1(46));
   U2684 : AOI221X2 port map( IN1 => RAM_12_46_port, IN2 => n2457, IN3 => 
                           RAM_13_46_port, IN4 => n3371, IN5 => n3012, QN => 
                           n2425);
   U2685 : AOI221X1 port map( IN1 => RAM_0_46_port, IN2 => n2170, IN3 => 
                           RAM_1_46_port, IN4 => n3384, IN5 => n3013, QN => 
                           n2426);
   U2686 : AOI221X2 port map( IN1 => RAM_4_46_port, IN2 => n3410, IN3 => 
                           RAM_5_46_port, IN4 => n3393, IN5 => n3014, QN => 
                           n2427);
   U2687 : AOI221X1 port map( IN1 => RAM_8_79_port, IN2 => n3424, IN3 => 
                           RAM_9_79_port, IN4 => n2493, IN5 => n3143, QN => 
                           n2672);
   U2688 : NAND4X0 port map( IN1 => n2428, IN2 => n2429, IN3 => n2430, IN4 => 
                           n2431, QN => RAMDOUT1(82));
   U2689 : AOI221X2 port map( IN1 => RAM_12_82_port, IN2 => n2450, IN3 => 
                           RAM_13_82_port, IN4 => n2490, IN5 => n3156, QN => 
                           n2429);
   U2690 : AOI221X1 port map( IN1 => RAM_0_82_port, IN2 => n2167, IN3 => 
                           RAM_1_82_port, IN4 => n3390, IN5 => n3157, QN => 
                           n2430);
   U2691 : AOI221X2 port map( IN1 => RAM_4_82_port, IN2 => n3448, IN3 => 
                           RAM_5_82_port, IN4 => n3400, IN5 => n3158, QN => 
                           n2431);
   U2692 : AO22X2 port map( IN1 => RAM_3_29_port, IN2 => n2550, IN3 => 
                           RAM_2_29_port, IN4 => n2643, Q => n2945);
   U2693 : AO22X2 port map( IN1 => RAM_3_112_port, IN2 => n2550, IN3 => 
                           RAM_2_112_port, IN4 => n2625, Q => n3277);
   U2694 : AO22X2 port map( IN1 => RAM_3_116_port, IN2 => n2542, IN3 => n2633, 
                           IN4 => RAM_2_116_port, Q => n3297);
   U2695 : AO22X2 port map( IN1 => RAM_3_46_port, IN2 => n2539, IN3 => n2640, 
                           IN4 => RAM_2_46_port, Q => n3013);
   U2696 : AO22X2 port map( IN1 => RAM_3_108_port, IN2 => n2538, IN3 => 
                           RAM_2_108_port, IN4 => n2111, Q => n3261);
   U2697 : AO22X2 port map( IN1 => RAM_3_125_port, IN2 => n2551, IN3 => 
                           RAM_2_125_port, IN4 => n2640, Q => n3333);
   U2698 : NAND4X0 port map( IN1 => n2432, IN2 => n2433, IN3 => n2434, IN4 => 
                           n2435, QN => RAMDOUT1(87));
   U2699 : AOI221X2 port map( IN1 => RAM_12_87_port, IN2 => n2446, IN3 => 
                           RAM_13_87_port, IN4 => n3380, IN5 => n3176, QN => 
                           n2433);
   U2700 : AOI221X2 port map( IN1 => RAM_4_87_port, IN2 => n3407, IN3 => 
                           RAM_5_87_port, IN4 => n2495, IN5 => n3178, QN => 
                           n2435);
   U2701 : NAND4X0 port map( IN1 => n2436, IN2 => n2437, IN3 => n2438, IN4 => 
                           n2439, QN => RAMDOUT1(109));
   U2702 : AOI221X2 port map( IN1 => RAM_12_109_port, IN2 => n2450, IN3 => 
                           RAM_13_109_port, IN4 => n3381, IN5 => n3264, QN => 
                           n2437);
   U2703 : AOI221X2 port map( IN1 => RAM_4_109_port, IN2 => n3405, IN3 => 
                           RAM_5_109_port, IN4 => n3391, IN5 => n3266, QN => 
                           n2439);
   U2704 : NAND4X0 port map( IN1 => n2440, IN2 => n2442, IN3 => n2441, IN4 => 
                           n2443, QN => RAMDOUT1(28));
   U2705 : AOI221X2 port map( IN1 => RAM_12_28_port, IN2 => n2460, IN3 => 
                           RAM_13_28_port, IN4 => n3373, IN5 => n2940, QN => 
                           n2441);
   U2706 : AOI221X1 port map( IN1 => RAM_0_28_port, IN2 => n2158, IN3 => 
                           RAM_1_28_port, IN4 => n3389, IN5 => n2941, QN => 
                           n2442);
   U2707 : AOI221X2 port map( IN1 => RAM_4_28_port, IN2 => n3408, IN3 => 
                           RAM_5_28_port, IN4 => n3398, IN5 => n2942, QN => 
                           n2443);
   U2708 : AO22X2 port map( IN1 => RAM_11_96_port, IN2 => n2504, IN3 => n2650, 
                           IN4 => RAM_10_96_port, Q => n3211);
   U2709 : AO22X2 port map( IN1 => RAM_11_106_port, IN2 => n2466, IN3 => 
                           RAM_10_106_port, IN4 => n2480, Q => n3251);
   U2710 : AND2X4 port map( IN1 => n2825, IN2 => n2821, Q => n2444);
   U2711 : NBUFFX2 port map( INP => n2444, Z => n2445);
   U2712 : NBUFFX2 port map( INP => n2444, Z => n2446);
   U2713 : NBUFFX2 port map( INP => n2444, Z => n2447);
   U2714 : NBUFFX2 port map( INP => n2444, Z => n2448);
   U2715 : NBUFFX2 port map( INP => n2444, Z => n2449);
   U2716 : NBUFFX2 port map( INP => n2444, Z => n2450);
   U2717 : NBUFFX2 port map( INP => n2444, Z => n2451);
   U2718 : NBUFFX2 port map( INP => n2444, Z => n2452);
   U2719 : DELLN1X2 port map( INP => n3347, Z => n2453);
   U2720 : DELLN1X2 port map( INP => n3347, Z => n2455);
   U2721 : DELLN1X2 port map( INP => n3347, Z => n2456);
   U2722 : NBUFFX2 port map( INP => n3347, Z => n2457);
   U2723 : DELLN1X2 port map( INP => n3347, Z => n2458);
   U2724 : DELLN1X2 port map( INP => n3347, Z => n2459);
   U2725 : INVX0 port map( INP => n3339, ZN => n2647);
   U2726 : INVX0 port map( INP => n2646, ZN => n2461);
   U2727 : INVX0 port map( INP => n3339, ZN => n2648);
   U2728 : INVX0 port map( INP => n2533, ZN => n2500);
   U2729 : NAND4X0 port map( IN1 => n2462, IN2 => n2463, IN3 => n2464, IN4 => 
                           n2465, QN => RAMDOUT1(47));
   U2730 : AOI221X2 port map( IN1 => RAM_12_47_port, IN2 => n2445, IN3 => 
                           RAM_13_47_port, IN4 => n3372, IN5 => n3016, QN => 
                           n2463);
   U2731 : AOI221X1 port map( IN1 => RAM_0_47_port, IN2 => n2158, IN3 => 
                           RAM_1_47_port, IN4 => n3386, IN5 => n3017, QN => 
                           n2464);
   U2732 : AOI221X2 port map( IN1 => RAM_4_47_port, IN2 => n3405, IN3 => 
                           RAM_5_47_port, IN4 => n3397, IN5 => n3018, QN => 
                           n2465);
   U2733 : INVX0 port map( INP => n3464, ZN => n2466);
   U2734 : INVX0 port map( INP => n3354, ZN => n2510);
   U2735 : INVX0 port map( INP => n2647, ZN => n2467);
   U2736 : INVX0 port map( INP => n2508, ZN => n2468);
   U2737 : INVX0 port map( INP => n3354, ZN => n2512);
   U2738 : INVX0 port map( INP => n2532, ZN => n2469);
   U2739 : INVX0 port map( INP => n3349, ZN => n2534);
   U2740 : INVX0 port map( INP => n2533, ZN => n2470);
   U2741 : INVX0 port map( INP => n3349, ZN => n2535);
   U2742 : NAND4X0 port map( IN1 => n2471, IN2 => n2472, IN3 => n2473, IN4 => 
                           n2474, QN => RAMDOUT1(80));
   U2743 : AOI221X2 port map( IN1 => RAM_12_80_port, IN2 => n2454, IN3 => 
                           RAM_13_80_port, IN4 => n2489, IN5 => n3148, QN => 
                           n2472);
   U2744 : AOI221X1 port map( IN1 => RAM_0_80_port, IN2 => n2161, IN3 => 
                           RAM_1_80_port, IN4 => n3386, IN5 => n3149, QN => 
                           n2473);
   U2745 : AOI221X2 port map( IN1 => RAM_4_80_port, IN2 => n3405, IN3 => 
                           RAM_5_80_port, IN4 => n3391, IN5 => n3150, QN => 
                           n2474);
   U2746 : NAND4X0 port map( IN1 => n2475, IN2 => n2476, IN3 => n2477, IN4 => 
                           n2478, QN => RAMDOUT1(63));
   U2747 : AOI221X2 port map( IN1 => RAM_12_63_port, IN2 => n2446, IN3 => 
                           RAM_13_63_port, IN4 => n3378, IN5 => n3080, QN => 
                           n2476);
   U2748 : AOI221X2 port map( IN1 => RAM_4_63_port, IN2 => n3403, IN3 => 
                           RAM_5_63_port, IN4 => n3397, IN5 => n3082, QN => 
                           n2478);
   U2749 : INVX0 port map( INP => n2535, ZN => n2479);
   U2750 : AO22X2 port map( IN1 => RAM_3_87_port, IN2 => n2549, IN3 => n2642, 
                           IN4 => RAM_2_87_port, Q => n3177);
   U2751 : INVX0 port map( INP => n2649, ZN => n2480);
   U2752 : INVX0 port map( INP => n3339, ZN => n2649);
   U2753 : INVX0 port map( INP => n2508, ZN => n2514);
   U2754 : INVX0 port map( INP => n2508, ZN => n2513);
   U2755 : NAND4X0 port map( IN1 => n2481, IN2 => n2482, IN3 => n2483, IN4 => 
                           n2484, QN => RAMDOUT1(122));
   U2756 : AOI221X2 port map( IN1 => RAM_12_122_port, IN2 => n2451, IN3 => 
                           RAM_13_122_port, IN4 => n2489, IN5 => n3320, QN => 
                           n2482);
   U2757 : AOI221X2 port map( IN1 => RAM_4_122_port, IN2 => n3403, IN3 => 
                           RAM_5_122_port, IN4 => n3397, IN5 => n3322, QN => 
                           n2484);
   U2758 : NAND4X0 port map( IN1 => n2485, IN2 => n2486, IN3 => n2487, IN4 => 
                           n2488, QN => RAMDOUT1(106));
   U2759 : AOI221X1 port map( IN1 => RAM_12_106_port, IN2 => n2456, IN3 => 
                           RAM_13_106_port, IN4 => n3376, IN5 => n3252, QN => 
                           n2486);
   U2760 : AOI221X1 port map( IN1 => RAM_0_106_port, IN2 => n2170, IN3 => 
                           RAM_1_106_port, IN4 => n2157, IN5 => n3253, QN => 
                           n2487);
   U2761 : AOI221X2 port map( IN1 => RAM_4_106_port, IN2 => n3403, IN3 => 
                           RAM_5_106_port, IN4 => n3399, IN5 => n3254, QN => 
                           n2488);
   U2762 : DELLN1X2 port map( INP => n3346, Z => n2489);
   U2763 : DELLN1X2 port map( INP => n3346, Z => n2490);
   U2764 : DELLN1X2 port map( INP => n3351, Z => n2491);
   U2765 : DELLN1X2 port map( INP => n3351, Z => n2492);
   U2766 : DELLN1X2 port map( INP => n3342, Z => n2493);
   U2767 : DELLN1X2 port map( INP => n3356, Z => n2494);
   U2768 : DELLN1X2 port map( INP => n3356, Z => n2495);
   U2769 : INVX0 port map( INP => n2647, ZN => n2653);
   U2770 : INVX0 port map( INP => n2648, ZN => n2651);
   U2771 : INVX0 port map( INP => n2649, ZN => n2652);
   U2772 : AO22X2 port map( IN1 => RAM_3_122_port, IN2 => n2554, IN3 => 
                           RAM_2_122_port, IN4 => n2623, Q => n3321);
   U2773 : AO22X2 port map( IN1 => RAM_3_95_port, IN2 => n2552, IN3 => 
                           RAM_2_95_port, IN4 => n2623, Q => n3209);
   U2774 : AO22X2 port map( IN1 => RAM_3_22_port, IN2 => n2546, IN3 => 
                           RAM_2_22_port, IN4 => n2643, Q => n2917);
   U2775 : AO22X2 port map( IN1 => RAM_3_44_port, IN2 => n2552, IN3 => 
                           RAM_2_44_port, IN4 => n2099, Q => n3005);
   U2776 : AOI221X1 port map( IN1 => RAM_0_22_port, IN2 => n2172, IN3 => 
                           RAM_1_22_port, IN4 => n2157, IN5 => n2917, QN => 
                           n2616);
   U2777 : AOI221X1 port map( IN1 => RAM_0_14_port, IN2 => n2160, IN3 => 
                           RAM_1_14_port, IN4 => n2492, IN5 => n2885, QN => 
                           n2580);
   U2778 : AOI221X1 port map( IN1 => RAM_0_13_port, IN2 => n2158, IN3 => 
                           RAM_1_13_port, IN4 => n2157, IN5 => n2881, QN => 
                           n2694);
   U2779 : AO22X2 port map( IN1 => RAM_3_63_port, IN2 => n2547, IN3 => 
                           RAM_2_63_port, IN4 => n2627, Q => n3081);
   U2780 : AO22X2 port map( IN1 => RAM_3_64_port, IN2 => n2547, IN3 => n2111, 
                           IN4 => RAM_2_64_port, Q => n3085);
   U2781 : AO22X2 port map( IN1 => RAM_3_119_port, IN2 => n2470, IN3 => n2111, 
                           IN4 => RAM_2_119_port, Q => n3309);
   U2782 : AO22X2 port map( IN1 => RAM_3_80_port, IN2 => n2545, IN3 => n2628, 
                           IN4 => RAM_2_80_port, Q => n3149);
   U2783 : AO22X2 port map( IN1 => RAM_3_110_port, IN2 => n2553, IN3 => n2628, 
                           IN4 => RAM_2_110_port, Q => n3269);
   U2784 : AO22X2 port map( IN1 => RAM_3_42_port, IN2 => n2470, IN3 => 
                           RAM_2_42_port, IN4 => n2624, Q => n2997);
   U2785 : AO22X2 port map( IN1 => RAM_3_32_port, IN2 => n2549, IN3 => 
                           RAM_2_32_port, IN4 => n2624, Q => n2957);
   U2786 : AO22X2 port map( IN1 => RAM_3_65_port, IN2 => n2546, IN3 => 
                           RAM_2_65_port, IN4 => n2630, Q => n3089);
   U2787 : AO22X2 port map( IN1 => RAM_3_61_port, IN2 => n2550, IN3 => 
                           RAM_2_61_port, IN4 => n2642, Q => n3073);
   U2788 : AO22X2 port map( IN1 => RAM_3_50_port, IN2 => n2540, IN3 => 
                           RAM_2_50_port, IN4 => n2632, Q => n3029);
   U2789 : AO22X2 port map( IN1 => RAM_3_104_port, IN2 => n2479, IN3 => 
                           RAM_2_104_port, IN4 => n2630, Q => n3245);
   U2790 : AO22X2 port map( IN1 => RAM_3_16_port, IN2 => n2500, IN3 => 
                           RAM_2_16_port, IN4 => n2625, Q => n2893);
   U2791 : AO22X2 port map( IN1 => RAM_3_126_port, IN2 => n2541, IN3 => 
                           RAM_2_126_port, IN4 => n2628, Q => n3337);
   U2792 : AO22X2 port map( IN1 => RAM_3_54_port, IN2 => n2544, IN3 => 
                           RAM_2_54_port, IN4 => n2634, Q => n3045);
   U2793 : AO22X2 port map( IN1 => RAM_3_67_port, IN2 => n2546, IN3 => 
                           RAM_2_67_port, IN4 => n2634, Q => n3097);
   U2794 : AO22X2 port map( IN1 => RAM_3_68_port, IN2 => n2543, IN3 => 
                           RAM_2_68_port, IN4 => n2639, Q => n3101);
   U2795 : AO22X2 port map( IN1 => RAM_3_33_port, IN2 => n2469, IN3 => 
                           RAM_2_33_port, IN4 => n2635, Q => n2961);
   U2796 : AO22X2 port map( IN1 => RAM_3_55_port, IN2 => n2540, IN3 => 
                           RAM_2_55_port, IN4 => n2635, Q => n3049);
   U2797 : AO22X2 port map( IN1 => RAM_3_107_port, IN2 => n2537, IN3 => 
                           RAM_2_107_port, IN4 => n2635, Q => n3257);
   U2798 : IBUFFX16 port map( INP => RAMADDR1(1), ZN => n2496);
   U2799 : INVX0 port map( INP => n2496, ZN => n2497);
   U2800 : AND2X4 port map( IN1 => n3359, IN2 => RAMADDR1(1), Q => n2797);
   U2801 : INVX0 port map( INP => n3463, ZN => n2498);
   U2802 : INVX0 port map( INP => n3340, ZN => n2499);
   U2803 : INVX0 port map( INP => n3349, ZN => n2533);
   U2804 : AND2X4 port map( IN1 => n2825, IN2 => n2819, Q => n3427);
   U2805 : INVX0 port map( INP => n2499, ZN => n2501);
   U2806 : NBUFFX2 port map( INP => RAMDIN1(99), Z => n2502);
   U2807 : NBUFFX2 port map( INP => RAMDIN1(99), Z => n2503);
   U2808 : AND2X1 port map( IN1 => n2823, IN2 => n2496, Q => n2505);
   U2809 : NBUFFX2 port map( INP => RAMDIN1(41), Z => n2506);
   U2810 : NBUFFX2 port map( INP => RAMDIN1(41), Z => n2507);
   U2811 : INVX0 port map( INP => n3354, ZN => n2508);
   U2812 : INVX0 port map( INP => n3354, ZN => n2509);
   U2813 : INVX0 port map( INP => n2508, ZN => n2515);
   U2814 : INVX0 port map( INP => n2508, ZN => n2516);
   U2815 : INVX0 port map( INP => n2509, ZN => n2517);
   U2816 : INVX0 port map( INP => n2509, ZN => n2518);
   U2817 : INVX0 port map( INP => n2509, ZN => n2519);
   U2818 : INVX0 port map( INP => n2509, ZN => n2520);
   U2819 : INVX0 port map( INP => n2510, ZN => n2521);
   U2820 : INVX0 port map( INP => n2510, ZN => n2522);
   U2821 : INVX0 port map( INP => n2510, ZN => n2523);
   U2822 : INVX0 port map( INP => n2510, ZN => n2524);
   U2823 : INVX0 port map( INP => n2511, ZN => n2525);
   U2824 : INVX0 port map( INP => n2511, ZN => n2526);
   U2825 : INVX0 port map( INP => n2511, ZN => n2527);
   U2826 : INVX0 port map( INP => n2512, ZN => n2528);
   U2827 : INVX0 port map( INP => n2512, ZN => n2529);
   U2828 : INVX0 port map( INP => n2512, ZN => n2530);
   U2829 : INVX0 port map( INP => n2512, ZN => n2531);
   U2830 : INVX0 port map( INP => n3349, ZN => n2532);
   U2831 : INVX0 port map( INP => n2532, ZN => n2538);
   U2832 : INVX0 port map( INP => n2535, ZN => n2539);
   U2833 : INVX0 port map( INP => n2536, ZN => n2540);
   U2834 : INVX0 port map( INP => n2533, ZN => n2541);
   U2835 : INVX0 port map( INP => n2536, ZN => n2542);
   U2836 : INVX0 port map( INP => n2535, ZN => n2543);
   U2837 : INVX0 port map( INP => n2536, ZN => n2544);
   U2838 : INVX0 port map( INP => n2535, ZN => n2545);
   U2839 : INVX0 port map( INP => n2532, ZN => n2546);
   U2840 : INVX0 port map( INP => n2534, ZN => n2547);
   U2841 : INVX0 port map( INP => n2533, ZN => n2548);
   U2842 : INVX0 port map( INP => n2535, ZN => n2549);
   U2843 : INVX0 port map( INP => n2536, ZN => n2550);
   U2844 : INVX0 port map( INP => n2534, ZN => n2551);
   U2845 : INVX0 port map( INP => n2532, ZN => n2552);
   U2846 : INVX0 port map( INP => n2533, ZN => n2553);
   U2847 : INVX0 port map( INP => n2534, ZN => n2554);
   U2848 : NBUFFX2 port map( INP => RAMDIN1(52), Z => n2555);
   U2849 : NBUFFX2 port map( INP => RAMDIN1(52), Z => n2556);
   U2850 : NBUFFX2 port map( INP => RAMDIN1(48), Z => n2557);
   U2851 : NBUFFX2 port map( INP => RAMDIN1(37), Z => n2558);
   U2852 : NBUFFX2 port map( INP => RAMDIN1(37), Z => n2559);
   U2853 : NBUFFX2 port map( INP => RAMDIN1(43), Z => n2560);
   U2854 : NBUFFX2 port map( INP => RAMDIN1(43), Z => n2561);
   U2855 : AOI221X2 port map( IN1 => RAM_12_59_port, IN2 => n2459, IN3 => 
                           RAM_13_59_port, IN4 => n3380, IN5 => n3064, QN => 
                           n2701);
   U2856 : DELLN1X2 port map( INP => n3346, Z => n3371);
   U2857 : DELLN1X2 port map( INP => n3346, Z => n3372);
   U2858 : DELLN1X2 port map( INP => n3346, Z => n3377);
   U2859 : DELLN1X2 port map( INP => n3346, Z => n3374);
   U2860 : DELLN1X2 port map( INP => n3346, Z => n3375);
   U2861 : DELLN1X2 port map( INP => n3346, Z => n3380);
   U2862 : NAND4X0 port map( IN1 => n2562, IN2 => n2563, IN3 => n2564, IN4 => 
                           n2565, QN => RAMDOUT1(42));
   U2863 : AOI221X2 port map( IN1 => RAM_12_42_port, IN2 => n2452, IN3 => 
                           RAM_13_42_port, IN4 => n3372, IN5 => n2996, QN => 
                           n2563);
   U2864 : AOI221X2 port map( IN1 => RAM_4_42_port, IN2 => n3405, IN3 => 
                           RAM_5_42_port, IN4 => n3395, IN5 => n2998, QN => 
                           n2565);
   U2865 : DELLN1X2 port map( INP => n3342, Z => n3360);
   U2866 : DELLN1X2 port map( INP => n3342, Z => n3363);
   U2867 : DELLN1X2 port map( INP => n3342, Z => n3364);
   U2868 : INVX0 port map( INP => n3339, ZN => n2646);
   U2869 : DELLN1X2 port map( INP => n3356, Z => n3391);
   U2870 : DELLN1X2 port map( INP => n3356, Z => n3394);
   U2871 : DELLN1X2 port map( INP => n3356, Z => n3393);
   U2872 : DELLN1X2 port map( INP => n3356, Z => n3401);
   U2873 : DELLN1X2 port map( INP => n3356, Z => n3399);
   U2874 : DELLN1X2 port map( INP => n3356, Z => n3395);
   U2875 : NAND4X0 port map( IN1 => n2566, IN2 => n2567, IN3 => n2568, IN4 => 
                           n2569, QN => RAMDOUT1(34));
   U2876 : AOI221X2 port map( IN1 => RAM_12_34_port, IN2 => n2458, IN3 => 
                           RAM_13_34_port, IN4 => n3375, IN5 => n2964, QN => 
                           n2567);
   U2877 : AOI221X2 port map( IN1 => RAM_4_34_port, IN2 => n3448, IN3 => 
                           RAM_5_34_port, IN4 => n3395, IN5 => n2966, QN => 
                           n2569);
   U2878 : NAND4X0 port map( IN1 => n2570, IN2 => n2571, IN3 => n2572, IN4 => 
                           n2573, QN => RAMDOUT1(39));
   U2879 : AOI221X2 port map( IN1 => RAM_12_39_port, IN2 => n2447, IN3 => 
                           RAM_13_39_port, IN4 => n3378, IN5 => n2984, QN => 
                           n2571);
   U2880 : AOI221X2 port map( IN1 => RAM_4_39_port, IN2 => n3407, IN3 => 
                           RAM_5_39_port, IN4 => n3393, IN5 => n2986, QN => 
                           n2573);
   U2881 : NAND4X0 port map( IN1 => n2574, IN2 => n2575, IN3 => n2576, IN4 => 
                           n2577, QN => RAMDOUT1(20));
   U2882 : AOI221X2 port map( IN1 => RAM_12_20_port, IN2 => n2451, IN3 => 
                           RAM_13_20_port, IN4 => n3374, IN5 => n2908, QN => 
                           n2575);
   U2883 : AOI221X2 port map( IN1 => RAM_4_20_port, IN2 => n3404, IN3 => 
                           RAM_5_20_port, IN4 => n3392, IN5 => n2910, QN => 
                           n2577);
   U2884 : NAND4X0 port map( IN1 => n2578, IN2 => n2579, IN3 => n2580, IN4 => 
                           n2581, QN => RAMDOUT1(14));
   U2885 : AOI221X2 port map( IN1 => RAM_12_14_port, IN2 => n2449, IN3 => 
                           RAM_13_14_port, IN4 => n3371, IN5 => n2884, QN => 
                           n2579);
   U2886 : AOI221X2 port map( IN1 => RAM_4_14_port, IN2 => n3408, IN3 => 
                           RAM_5_14_port, IN4 => n3396, IN5 => n2886, QN => 
                           n2581);
   U2887 : DELLN1X2 port map( INP => n3351, Z => n3382);
   U2888 : DELLN1X2 port map( INP => n3351, Z => n3389);
   U2889 : DELLN1X2 port map( INP => n3351, Z => n3390);
   U2890 : DELLN1X2 port map( INP => n3351, Z => n3385);
   U2891 : NAND4X0 port map( IN1 => n2582, IN2 => n2583, IN3 => n2584, IN4 => 
                           n2585, QN => RAMDOUT1(38));
   U2892 : AOI221X2 port map( IN1 => RAM_12_38_port, IN2 => n2460, IN3 => 
                           RAM_13_38_port, IN4 => n3380, IN5 => n2980, QN => 
                           n2583);
   U2893 : AOI221X2 port map( IN1 => RAM_4_38_port, IN2 => n3407, IN3 => 
                           RAM_5_38_port, IN4 => n3395, IN5 => n2982, QN => 
                           n2585);
   U2894 : NAND4X0 port map( IN1 => n2586, IN2 => n2587, IN3 => n2588, IN4 => 
                           n2589, QN => RAMDOUT1(45));
   U2895 : AOI221X2 port map( IN1 => RAM_12_45_port, IN2 => n2446, IN3 => 
                           RAM_13_45_port, IN4 => n3373, IN5 => n3008, QN => 
                           n2587);
   U2896 : AOI221X2 port map( IN1 => RAM_4_45_port, IN2 => n3409, IN3 => 
                           RAM_5_45_port, IN4 => n3399, IN5 => n3010, QN => 
                           n2589);
   U2897 : AO22X2 port map( IN1 => RAM_15_96_port, IN2 => n3435, IN3 => 
                           RAM_14_96_port, IN4 => n2322, Q => n3212);
   U2898 : NAND4X0 port map( IN1 => n2590, IN2 => n2591, IN3 => n2592, IN4 => 
                           n2593, QN => RAMDOUT1(4));
   U2899 : AOI221X2 port map( IN1 => RAM_12_4_port, IN2 => n2455, IN3 => 
                           RAM_13_4_port, IN4 => n3377, IN5 => n2844, QN => 
                           n2591);
   U2900 : AOI221X2 port map( IN1 => RAM_4_4_port, IN2 => n3404, IN3 => 
                           RAM_5_4_port, IN4 => n3399, IN5 => n2846, QN => 
                           n2593);
   U2901 : NAND4X0 port map( IN1 => n2594, IN2 => n2595, IN3 => n2596, IN4 => 
                           n2597, QN => RAMDOUT1(114));
   U2902 : AOI221X2 port map( IN1 => RAM_12_114_port, IN2 => n2457, IN3 => 
                           RAM_13_114_port, IN4 => n3381, IN5 => n3288, QN => 
                           n2595);
   U2903 : AOI221X2 port map( IN1 => RAM_4_114_port, IN2 => n3402, IN3 => 
                           RAM_5_114_port, IN4 => n3392, IN5 => n3290, QN => 
                           n2597);
   U2904 : AO22X2 port map( IN1 => RAM_15_109_port, IN2 => n3439, IN3 => 
                           RAM_14_109_port, IN4 => n2327, Q => n3264);
   U2905 : INVX0 port map( INP => n2618, ZN => n2631);
   U2906 : NAND4X0 port map( IN1 => n2598, IN2 => n2599, IN3 => n2600, IN4 => 
                           n2601, QN => RAMDOUT1(118));
   U2907 : AOI221X2 port map( IN1 => RAM_12_118_port, IN2 => n2456, IN3 => 
                           RAM_13_118_port, IN4 => n3376, IN5 => n3304, QN => 
                           n2599);
   U2908 : AOI221X2 port map( IN1 => RAM_4_118_port, IN2 => n3405, IN3 => 
                           RAM_5_118_port, IN4 => n3396, IN5 => n3306, QN => 
                           n2601);
   U2909 : NAND4X0 port map( IN1 => n2602, IN2 => n2603, IN3 => n2604, IN4 => 
                           n2605, QN => RAMDOUT1(56));
   U2910 : AOI221X2 port map( IN1 => RAM_12_56_port, IN2 => n2458, IN3 => 
                           RAM_13_56_port, IN4 => n3381, IN5 => n3052, QN => 
                           n2603);
   U2911 : AOI221X2 port map( IN1 => RAM_4_56_port, IN2 => n3408, IN3 => 
                           RAM_5_56_port, IN4 => n3399, IN5 => n3054, QN => 
                           n2605);
   U2912 : NAND4X0 port map( IN1 => n2606, IN2 => n2607, IN3 => n2608, IN4 => 
                           n2609, QN => RAMDOUT1(49));
   U2913 : AOI221X2 port map( IN1 => RAM_12_49_port, IN2 => n2450, IN3 => 
                           RAM_13_49_port, IN4 => n2489, IN5 => n3024, QN => 
                           n2607);
   U2914 : AOI221X2 port map( IN1 => RAM_4_49_port, IN2 => n3402, IN3 => 
                           RAM_5_49_port, IN4 => n3400, IN5 => n3026, QN => 
                           n2609);
   U2915 : NAND4X0 port map( IN1 => n2610, IN2 => n2611, IN3 => n2612, IN4 => 
                           n2613, QN => RAMDOUT1(94));
   U2916 : AOI221X2 port map( IN1 => RAM_12_94_port, IN2 => n2450, IN3 => 
                           RAM_13_94_port, IN4 => n2490, IN5 => n3204, QN => 
                           n2612);
   U2917 : AOI221X2 port map( IN1 => RAM_4_94_port, IN2 => n3407, IN3 => 
                           RAM_5_94_port, IN4 => n3400, IN5 => n3206, QN => 
                           n2613);
   U2918 : DELLN1X2 port map( INP => n3346, Z => n3373);
   U2919 : AO22X2 port map( IN1 => RAM_15_34_port, IN2 => n3444, IN3 => 
                           RAM_14_34_port, IN4 => n2334, Q => n2964);
   U2920 : AO22X2 port map( IN1 => RAM_15_78_port, IN2 => n3433, IN3 => 
                           RAM_14_78_port, IN4 => n2336, Q => n3140);
   U2921 : AO22X2 port map( IN1 => RAM_15_7_port, IN2 => n3438, IN3 => 
                           RAM_14_7_port, IN4 => n2328, Q => n2856);
   U2922 : AO22X2 port map( IN1 => RAM_15_30_port, IN2 => n3444, IN3 => 
                           RAM_14_30_port, IN4 => n2331, Q => n2948);
   U2923 : OR4X2 port map( IN1 => n4240, IN2 => n4239, IN3 => n4238, IN4 => 
                           n4237, Q => RAMDOUT2(95));
   U2924 : AO22X2 port map( IN1 => RAM_15_81_port, IN2 => n3438, IN3 => 
                           RAM_14_81_port, IN4 => n2335, Q => n3152);
   U2925 : AO22X2 port map( IN1 => RAM_15_89_port, IN2 => n3445, IN3 => 
                           RAM_14_89_port, IN4 => n2326, Q => n3184);
   U2926 : AO22X2 port map( IN1 => RAM_15_47_port, IN2 => n3436, IN3 => 
                           RAM_14_47_port, IN4 => n2324, Q => n3016);
   U2927 : AO22X2 port map( IN1 => RAM_15_44_port, IN2 => n3440, IN3 => 
                           RAM_14_44_port, IN4 => n2331, Q => n3004);
   U2928 : AO22X2 port map( IN1 => RAM_15_57_port, IN2 => n3433, IN3 => 
                           RAM_14_57_port, IN4 => n2334, Q => n3056);
   U2929 : AO22X2 port map( IN1 => RAM_15_0_port, IN2 => n3444, IN3 => 
                           RAM_14_0_port, IN4 => n2334, Q => n2822);
   U2930 : NAND4X0 port map( IN1 => n2614, IN2 => n2615, IN3 => n2616, IN4 => 
                           n2617, QN => RAMDOUT1(22));
   U2931 : AOI221X1 port map( IN1 => RAM_8_22_port, IN2 => n3426, IN3 => 
                           RAM_9_22_port, IN4 => n3361, IN5 => n2915, QN => 
                           n2614);
   U2932 : AOI221X1 port map( IN1 => RAM_12_22_port, IN2 => n2446, IN3 => 
                           RAM_13_22_port, IN4 => n3379, IN5 => n2916, QN => 
                           n2615);
   U2933 : AOI221X1 port map( IN1 => RAM_4_22_port, IN2 => n3409, IN3 => 
                           RAM_5_22_port, IN4 => n3395, IN5 => n2918, QN => 
                           n2617);
   U2934 : AND2X4 port map( IN1 => n34, IN2 => n2708, Q => n25);
   U2935 : INVX0 port map( INP => n3348, ZN => n2618);
   U2936 : INVX0 port map( INP => n3348, ZN => n2619);
   U2937 : INVX0 port map( INP => n2622, ZN => n2623);
   U2938 : INVX0 port map( INP => n2618, ZN => n2624);
   U2939 : INVX0 port map( INP => n2620, ZN => n2625);
   U2940 : INVX0 port map( INP => n2621, ZN => n2626);
   U2941 : INVX0 port map( INP => n2621, ZN => n2627);
   U2942 : INVX0 port map( INP => n2619, ZN => n2628);
   U2943 : INVX0 port map( INP => n2618, ZN => n2629);
   U2944 : INVX0 port map( INP => n2620, ZN => n2630);
   U2945 : INVX0 port map( INP => n2620, ZN => n2632);
   U2946 : INVX0 port map( INP => n2619, ZN => n2633);
   U2947 : INVX0 port map( INP => n2622, ZN => n2635);
   U2948 : INVX0 port map( INP => n2618, ZN => n2636);
   U2949 : INVX0 port map( INP => n2622, ZN => n2637);
   U2950 : INVX0 port map( INP => n2621, ZN => n2639);
   U2951 : INVX0 port map( INP => n2621, ZN => n2640);
   U2952 : INVX0 port map( INP => n2619, ZN => n2641);
   U2953 : INVX0 port map( INP => n2620, ZN => n2642);
   U2954 : AO22X2 port map( IN1 => RAM_3_111_port, IN2 => n2399, IN3 => n2643, 
                           IN4 => RAM_2_111_port, Q => n3273);
   U2955 : AO22X2 port map( IN1 => RAM_3_106_port, IN2 => n2469, IN3 => n2623, 
                           IN4 => RAM_2_106_port, Q => n3253);
   U2956 : AO22X2 port map( IN1 => RAM_3_36_port, IN2 => n2538, IN3 => 
                           RAM_2_36_port, IN4 => n2639, Q => n2973);
   U2957 : AO22X2 port map( IN1 => RAM_3_17_port, IN2 => n2545, IN3 => 
                           RAM_2_17_port, IN4 => n2638, Q => n2897);
   U2958 : INVX0 port map( INP => n3339, ZN => n2645);
   U2959 : INVX0 port map( INP => n2649, ZN => n2650);
   U2960 : INVX0 port map( INP => n2646, ZN => n2655);
   U2961 : INVX0 port map( INP => n2649, ZN => n2656);
   U2962 : INVX0 port map( INP => n2645, ZN => n2657);
   U2963 : INVX0 port map( INP => n2648, ZN => n2658);
   U2964 : INVX0 port map( INP => n2648, ZN => n2659);
   U2965 : INVX0 port map( INP => n2647, ZN => n2660);
   U2966 : INVX0 port map( INP => n2645, ZN => n2661);
   U2967 : INVX0 port map( INP => n2645, ZN => n2662);
   U2968 : INVX0 port map( INP => n2648, ZN => n2664);
   U2969 : INVX0 port map( INP => n2646, ZN => n2665);
   U2970 : INVX0 port map( INP => n2648, ZN => n2667);
   U2971 : NAND4X0 port map( IN1 => n2668, IN2 => n2669, IN3 => n2670, IN4 => 
                           n2671, QN => RAMDOUT1(53));
   U2972 : AOI221X1 port map( IN1 => RAM_8_53_port, IN2 => n3417, IN3 => 
                           RAM_9_53_port, IN4 => n3365, IN5 => n3039, QN => 
                           n2668);
   U2973 : AOI221X2 port map( IN1 => RAM_12_53_port, IN2 => n2448, IN3 => 
                           RAM_13_53_port, IN4 => n3372, IN5 => n3040, QN => 
                           n2669);
   U2974 : AOI221X2 port map( IN1 => RAM_4_53_port, IN2 => n3405, IN3 => 
                           RAM_5_53_port, IN4 => n3392, IN5 => n3042, QN => 
                           n2671);
   U2975 : NAND4X0 port map( IN1 => n2672, IN2 => n2673, IN3 => n2674, IN4 => 
                           n2675, QN => RAMDOUT1(79));
   U2976 : AOI221X2 port map( IN1 => RAM_12_79_port, IN2 => n2459, IN3 => 
                           RAM_13_79_port, IN4 => n3374, IN5 => n3144, QN => 
                           n2673);
   U2977 : AOI221X2 port map( IN1 => RAM_4_79_port, IN2 => n3404, IN3 => 
                           RAM_5_79_port, IN4 => n2494, IN5 => n3146, QN => 
                           n2675);
   U2978 : NAND4X0 port map( IN1 => n2676, IN2 => n2677, IN3 => n2678, IN4 => 
                           n2679, QN => RAMDOUT1(78));
   U2979 : AOI221X2 port map( IN1 => RAM_12_78_port, IN2 => n2445, IN3 => 
                           RAM_13_78_port, IN4 => n3379, IN5 => n3140, QN => 
                           n2677);
   U2980 : AOI221X2 port map( IN1 => RAM_4_78_port, IN2 => n3448, IN3 => 
                           RAM_5_78_port, IN4 => n3391, IN5 => n3142, QN => 
                           n2679);
   U2981 : NAND4X0 port map( IN1 => n2680, IN2 => n2681, IN3 => n2682, IN4 => 
                           n2683, QN => RAMDOUT1(51));
   U2982 : AOI221X1 port map( IN1 => RAM_8_51_port, IN2 => n3420, IN3 => 
                           RAM_9_51_port, IN4 => n3363, IN5 => n3031, QN => 
                           n2680);
   U2983 : AOI221X1 port map( IN1 => RAM_0_51_port, IN2 => n2171, IN3 => 
                           RAM_1_51_port, IN4 => n3389, IN5 => n3033, QN => 
                           n2682);
   U2984 : AOI221X1 port map( IN1 => RAM_4_51_port, IN2 => n3402, IN3 => 
                           RAM_5_51_port, IN4 => n3400, IN5 => n3034, QN => 
                           n2683);
   U2985 : NAND4X0 port map( IN1 => n2686, IN2 => n2685, IN3 => n2684, IN4 => 
                           n2687, QN => RAMDOUT1(61));
   U2986 : AOI221X1 port map( IN1 => RAM_8_61_port, IN2 => n3415, IN3 => 
                           RAM_9_61_port, IN4 => n3361, IN5 => n3071, QN => 
                           n2684);
   U2987 : AOI221X1 port map( IN1 => RAM_12_61_port, IN2 => n2450, IN3 => 
                           RAM_13_61_port, IN4 => n3381, IN5 => n3072, QN => 
                           n2685);
   U2988 : AOI221X1 port map( IN1 => RAM_0_61_port, IN2 => n2164, IN3 => 
                           RAM_1_61_port, IN4 => n3388, IN5 => n3073, QN => 
                           n2686);
   U2989 : AOI221X1 port map( IN1 => RAM_4_61_port, IN2 => n3403, IN3 => 
                           RAM_5_61_port, IN4 => n3396, IN5 => n3074, QN => 
                           n2687);
   U2990 : NAND4X0 port map( IN1 => n2688, IN2 => n2689, IN3 => n2690, IN4 => 
                           n2691, QN => RAMDOUT1(0));
   U2991 : AOI221X1 port map( IN1 => RAM_8_0_port, IN2 => n3424, IN3 => 
                           RAM_9_0_port, IN4 => n3363, IN5 => n2820, QN => 
                           n2688);
   U2992 : AOI221X1 port map( IN1 => RAM_12_0_port, IN2 => n2448, IN3 => 
                           RAM_13_0_port, IN4 => n2489, IN5 => n2822, QN => 
                           n2689);
   U2993 : AOI221X1 port map( IN1 => RAM_0_0_port, IN2 => n2161, IN3 => 
                           RAM_1_0_port, IN4 => n3385, IN5 => n2824, QN => 
                           n2690);
   U2994 : AOI221X2 port map( IN1 => RAM_4_0_port, IN2 => n3406, IN3 => 
                           RAM_5_0_port, IN4 => n3400, IN5 => n2830, QN => 
                           n2691);
   U2995 : NAND4X0 port map( IN1 => n2692, IN2 => n2693, IN3 => n2694, IN4 => 
                           n2695, QN => RAMDOUT1(13));
   U2996 : AOI221X1 port map( IN1 => RAM_8_13_port, IN2 => n3426, IN3 => 
                           RAM_9_13_port, IN4 => n3366, IN5 => n2879, QN => 
                           n2692);
   U2997 : AOI221X1 port map( IN1 => RAM_12_13_port, IN2 => n2454, IN3 => 
                           RAM_13_13_port, IN4 => n3371, IN5 => n2880, QN => 
                           n2693);
   U2998 : AOI221X1 port map( IN1 => RAM_4_13_port, IN2 => n3448, IN3 => 
                           RAM_5_13_port, IN4 => n3397, IN5 => n2882, QN => 
                           n2695);
   U2999 : NAND4X0 port map( IN1 => n2696, IN2 => n2697, IN3 => n2698, IN4 => 
                           n2699, QN => RAMDOUT1(32));
   U3000 : AOI221X1 port map( IN1 => RAM_8_32_port, IN2 => n3426, IN3 => 
                           RAM_9_32_port, IN4 => n3365, IN5 => n2955, QN => 
                           n2696);
   U3001 : AOI221X1 port map( IN1 => RAM_12_32_port, IN2 => n2451, IN3 => 
                           RAM_13_32_port, IN4 => n3380, IN5 => n2956, QN => 
                           n2697);
   U3002 : AOI221X1 port map( IN1 => RAM_0_32_port, IN2 => n2158, IN3 => 
                           RAM_1_32_port, IN4 => n3389, IN5 => n2957, QN => 
                           n2698);
   U3003 : AOI221X1 port map( IN1 => RAM_4_32_port, IN2 => n3403, IN3 => 
                           RAM_5_32_port, IN4 => n3401, IN5 => n2958, QN => 
                           n2699);
   U3004 : NAND4X0 port map( IN1 => n2700, IN2 => n2701, IN3 => n2702, IN4 => 
                           n2703, QN => RAMDOUT1(59));
   U3005 : AOI221X1 port map( IN1 => RAM_0_59_port, IN2 => n2166, IN3 => 
                           RAM_1_59_port, IN4 => n3390, IN5 => n3065, QN => 
                           n2702);
   U3006 : AOI221X1 port map( IN1 => RAM_4_59_port, IN2 => n3410, IN3 => 
                           RAM_5_59_port, IN4 => n3392, IN5 => n3066, QN => 
                           n2703);
   U3007 : NAND4X0 port map( IN1 => n2704, IN2 => n2705, IN3 => n2706, IN4 => 
                           n2707, QN => RAMDOUT1(8));
   U3008 : AOI221X1 port map( IN1 => RAM_8_8_port, IN2 => n3421, IN3 => 
                           RAM_9_8_port, IN4 => n3365, IN5 => n2859, QN => 
                           n2704);
   U3009 : AOI221X1 port map( IN1 => RAM_12_8_port, IN2 => n2447, IN3 => 
                           RAM_13_8_port, IN4 => n3375, IN5 => n2860, QN => 
                           n2705);
   U3010 : AOI221X1 port map( IN1 => RAM_0_8_port, IN2 => n2159, IN3 => 
                           RAM_1_8_port, IN4 => n2492, IN5 => n2861, QN => 
                           n2706);
   U3011 : AOI221X1 port map( IN1 => RAM_4_8_port, IN2 => n3408, IN3 => 
                           RAM_5_8_port, IN4 => n3401, IN5 => n2862, QN => 
                           n2707);
   U3012 : AO22X2 port map( IN1 => RAM_11_50_port, IN2 => n2498, IN3 => n2656, 
                           IN4 => RAM_10_50_port, Q => n3027);
   U3013 : AO22X1 port map( IN1 => RAM_7_90_port, IN2 => n2524, IN3 => 
                           RAM_6_90_port, IN4 => n2138, Q => n3190);
   U3014 : AO22X1 port map( IN1 => RAM_7_86_port, IN2 => n2523, IN3 => 
                           RAM_6_86_port, IN4 => n2150, Q => n3174);
   U3015 : AO22X1 port map( IN1 => RAM_7_95_port, IN2 => n2394, IN3 => 
                           RAM_6_95_port, IN4 => n2145, Q => n3210);
   U3016 : INVX0 port map( INP => n2708, ZN => n2709);
   U3017 : AO22X2 port map( IN1 => RAM_11_35_port, IN2 => n3453, IN3 => 
                           RAM_10_35_port, IN4 => n2663, Q => n2967);
   U3018 : AO22X2 port map( IN1 => RAM_11_39_port, IN2 => n3455, IN3 => n2662, 
                           IN4 => RAM_10_39_port, Q => n2983);
   U3019 : NAND4X0 port map( IN1 => n2710, IN2 => n2711, IN3 => n2712, IN4 => 
                           n2713, QN => RAMDOUT1(107));
   U3020 : AOI221X2 port map( IN1 => RAM_12_107_port, IN2 => n2452, IN3 => 
                           RAM_13_107_port, IN4 => n3381, IN5 => n3256, QN => 
                           n2711);
   U3021 : AOI221X1 port map( IN1 => RAM_0_69_port, IN2 => n2165, IN3 => 
                           RAM_1_69_port, IN4 => n2491, IN5 => n3105, QN => 
                           n2728);
   U3022 : AO22X2 port map( IN1 => RAM_11_90_port, IN2 => n3460, IN3 => n2658, 
                           IN4 => RAM_10_90_port, Q => n3187);
   U3023 : AO22X2 port map( IN1 => RAM_3_49_port, IN2 => n2541, IN3 => 
                           RAM_2_49_port, IN4 => n2629, Q => n3025);
   U3024 : AO22X2 port map( IN1 => RAM_3_77_port, IN2 => n2537, IN3 => 
                           RAM_2_77_port, IN4 => n2634, Q => n3137);
   U3025 : AO22X2 port map( IN1 => RAM_3_127_port, IN2 => n2540, IN3 => n2644, 
                           IN4 => RAM_2_127_port, Q => n3350);
   U3026 : AO22X2 port map( IN1 => RAM_11_0_port, IN2 => n3450, IN3 => 
                           RAM_10_0_port, IN4 => n2657, Q => n2820);
   U3027 : AOI221X1 port map( IN1 => RAM_8_101_port, IN2 => n3418, IN3 => 
                           RAM_9_101_port, IN4 => n3364, IN5 => n3231, QN => 
                           n2734);
   U3028 : NAND4X0 port map( IN1 => n2714, IN2 => n2715, IN3 => n2716, IN4 => 
                           n2717, QN => RAMDOUT1(76));
   U3029 : AOI221X2 port map( IN1 => RAM_12_76_port, IN2 => n2453, IN3 => 
                           RAM_13_76_port, IN4 => n3374, IN5 => n3132, QN => 
                           n2715);
   U3030 : AOI221X2 port map( IN1 => RAM_4_76_port, IN2 => n3409, IN3 => 
                           RAM_5_76_port, IN4 => n3399, IN5 => n3134, QN => 
                           n2717);
   U3031 : AO22X2 port map( IN1 => RAM_3_99_port, IN2 => n2542, IN3 => 
                           RAM_2_99_port, IN4 => n2636, Q => n3225);
   U3032 : AO22X2 port map( IN1 => RAM_3_91_port, IN2 => n2547, IN3 => 
                           RAM_2_91_port, IN4 => n2630, Q => n3193);
   U3033 : DELLN1X2 port map( INP => n3351, Z => n3383);
   U3034 : AO22X2 port map( IN1 => RAM_3_75_port, IN2 => n2551, IN3 => n2111, 
                           IN4 => RAM_2_75_port, Q => n3129);
   U3035 : AO22X2 port map( IN1 => RAM_3_79_port, IN2 => n2542, IN3 => 
                           RAM_2_79_port, IN4 => n2635, Q => n3145);
   U3036 : AO22X2 port map( IN1 => RAM_3_82_port, IN2 => n2544, IN3 => 
                           RAM_2_82_port, IN4 => n2637, Q => n3157);
   U3037 : AO22X2 port map( IN1 => RAM_3_94_port, IN2 => n2554, IN3 => 
                           RAM_2_94_port, IN4 => n2625, Q => n3205);
   U3038 : NAND4X0 port map( IN1 => n2718, IN2 => n2719, IN3 => n2720, IN4 => 
                           n2721, QN => RAMDOUT1(124));
   U3039 : AOI221X1 port map( IN1 => RAM_8_124_port, IN2 => n3420, IN3 => 
                           RAM_9_124_port, IN4 => n2493, IN5 => n3327, QN => 
                           n2718);
   U3040 : AOI221X1 port map( IN1 => RAM_12_124_port, IN2 => n2457, IN3 => 
                           RAM_13_124_port, IN4 => n3379, IN5 => n3328, QN => 
                           n2719);
   U3041 : AOI221X1 port map( IN1 => RAM_0_124_port, IN2 => n2164, IN3 => 
                           RAM_1_124_port, IN4 => n3382, IN5 => n3329, QN => 
                           n2720);
   U3042 : NAND4X0 port map( IN1 => n2722, IN2 => n2723, IN3 => n2724, IN4 => 
                           n2725, QN => RAMDOUT1(84));
   U3043 : AOI221X1 port map( IN1 => RAM_8_84_port, IN2 => n3422, IN3 => 
                           RAM_9_84_port, IN4 => n3363, IN5 => n3163, QN => 
                           n2722);
   U3044 : AOI221X2 port map( IN1 => RAM_12_84_port, IN2 => n2453, IN3 => 
                           RAM_13_84_port, IN4 => n2489, IN5 => n3164, QN => 
                           n2723);
   U3045 : AOI221X2 port map( IN1 => RAM_4_84_port, IN2 => n3408, IN3 => 
                           RAM_5_84_port, IN4 => n2495, IN5 => n3166, QN => 
                           n2725);
   U3046 : NAND4X0 port map( IN1 => n2726, IN2 => n2727, IN3 => n2728, IN4 => 
                           n2729, QN => RAMDOUT1(69));
   U3047 : AOI221X2 port map( IN1 => RAM_12_69_port, IN2 => n2460, IN3 => 
                           RAM_13_69_port, IN4 => n3373, IN5 => n3104, QN => 
                           n2727);
   U3048 : AOI221X2 port map( IN1 => RAM_4_69_port, IN2 => n3402, IN3 => 
                           RAM_5_69_port, IN4 => n3394, IN5 => n3106, QN => 
                           n2729);
   U3049 : NAND4X0 port map( IN1 => n2730, IN2 => n2731, IN3 => n2732, IN4 => 
                           n2733, QN => RAMDOUT1(25));
   U3050 : AOI221X2 port map( IN1 => RAM_8_25_port, IN2 => n3426, IN3 => 
                           RAM_9_25_port, IN4 => n3362, IN5 => n2927, QN => 
                           n2730);
   U3051 : AOI221X2 port map( IN1 => RAM_12_25_port, IN2 => n2455, IN3 => 
                           RAM_13_25_port, IN4 => n3377, IN5 => n2928, QN => 
                           n2731);
   U3052 : AOI221X1 port map( IN1 => RAM_0_25_port, IN2 => n2162, IN3 => 
                           RAM_1_25_port, IN4 => n2491, IN5 => n2929, QN => 
                           n2732);
   U3053 : AOI221X2 port map( IN1 => RAM_4_25_port, IN2 => n3448, IN3 => 
                           RAM_5_25_port, IN4 => n2495, IN5 => n2930, QN => 
                           n2733);
   U3054 : AO22X2 port map( IN1 => RAM_3_89_port, IN2 => n2539, IN3 => 
                           RAM_2_89_port, IN4 => n2626, Q => n3185);
   U3055 : AO22X2 port map( IN1 => RAM_3_84_port, IN2 => n2469, IN3 => n2641, 
                           IN4 => RAM_2_84_port, Q => n3165);
   U3056 : AO22X2 port map( IN1 => RAM_3_72_port, IN2 => n2399, IN3 => 
                           RAM_2_72_port, IN4 => n2642, Q => n3117);
   U3057 : AO22X2 port map( IN1 => RAM_3_31_port, IN2 => n2470, IN3 => 
                           RAM_2_31_port, IN4 => n2641, Q => n2953);
   U3058 : NAND4X0 port map( IN1 => n2734, IN2 => n2735, IN3 => n2737, IN4 => 
                           n2736, QN => RAMDOUT1(101));
   U3059 : AOI221X2 port map( IN1 => RAM_12_101_port, IN2 => n2450, IN3 => 
                           RAM_13_101_port, IN4 => n2489, IN5 => n3232, QN => 
                           n2735);
   U3060 : AOI221X2 port map( IN1 => RAM_4_101_port, IN2 => n3406, IN3 => 
                           RAM_5_101_port, IN4 => n3392, IN5 => n3234, QN => 
                           n2737);
   U3061 : AO22X2 port map( IN1 => RAM_3_34_port, IN2 => n2543, IN3 => n2641, 
                           IN4 => RAM_2_34_port, Q => n2965);
   U3062 : AO22X2 port map( IN1 => RAM_3_3_port, IN2 => n2549, IN3 => 
                           RAM_2_3_port, IN4 => n2626, Q => n2841);
   U3063 : AO22X2 port map( IN1 => RAM_3_13_port, IN2 => n2537, IN3 => 
                           RAM_2_13_port, IN4 => n2642, Q => n2881);
   U3064 : AO22X2 port map( IN1 => RAM_3_120_port, IN2 => n2554, IN3 => 
                           RAM_2_120_port, IN4 => n2625, Q => n3313);
   U3065 : AO22X2 port map( IN1 => RAM_3_43_port, IN2 => n2544, IN3 => 
                           RAM_2_43_port, IN4 => n2644, Q => n3001);
   U3066 : AO22X2 port map( IN1 => RAM_3_121_port, IN2 => n2539, IN3 => 
                           RAM_2_121_port, IN4 => n2632, Q => n3317);
   U3067 : AO22X2 port map( IN1 => RAM_3_60_port, IN2 => n2479, IN3 => 
                           RAM_2_60_port, IN4 => n2640, Q => n3069);
   U3068 : AO22X2 port map( IN1 => RAM_3_8_port, IN2 => n2553, IN3 => n2633, 
                           IN4 => RAM_2_8_port, Q => n2861);
   U3069 : AO22X2 port map( IN1 => RAM_3_100_port, IN2 => n2479, IN3 => n2629, 
                           IN4 => RAM_2_100_port, Q => n3229);
   U3070 : AO22X2 port map( IN1 => RAM_3_26_port, IN2 => n2553, IN3 => 
                           RAM_2_26_port, IN4 => n2624, Q => n2933);
   U3071 : NAND4X0 port map( IN1 => n2738, IN2 => n2739, IN3 => n2740, IN4 => 
                           n2741, QN => RAMDOUT1(126));
   U3072 : AOI221X1 port map( IN1 => RAM_8_126_port, IN2 => n3421, IN3 => 
                           RAM_9_126_port, IN4 => n3365, IN5 => n3335, QN => 
                           n2738);
   U3073 : AOI221X1 port map( IN1 => RAM_0_126_port, IN2 => n2163, IN3 => 
                           RAM_1_126_port, IN4 => n2491, IN5 => n3337, QN => 
                           n2740);
   U3074 : AOI221X1 port map( IN1 => RAM_4_126_port, IN2 => n3405, IN3 => 
                           RAM_5_126_port, IN4 => n3393, IN5 => n3338, QN => 
                           n2741);
   U3075 : AO22X2 port map( IN1 => RAM_3_69_port, IN2 => n2537, IN3 => 
                           RAM_2_69_port, IN4 => n2639, Q => n3105);
   U3076 : AO22X2 port map( IN1 => RAM_11_91_port, IN2 => n3453, IN3 => 
                           RAM_10_91_port, IN4 => n2652, Q => n3191);
   U3077 : AO22X2 port map( IN1 => RAM_3_117_port, IN2 => n2548, IN3 => 
                           RAM_2_117_port, IN4 => n2638, Q => n3301);
   U3078 : AO22X2 port map( IN1 => RAM_3_15_port, IN2 => n2542, IN3 => 
                           RAM_2_15_port, IN4 => n2634, Q => n2889);
   U3079 : AO22X2 port map( IN1 => RAM_3_86_port, IN2 => n2540, IN3 => 
                           RAM_2_86_port, IN4 => n2636, Q => n3173);
   U3080 : AO22X2 port map( IN1 => RAM_3_124_port, IN2 => n2552, IN3 => n2628, 
                           IN4 => RAM_2_124_port, Q => n3329);
   U3081 : AO22X2 port map( IN1 => RAM_3_59_port, IN2 => n2539, IN3 => 
                           RAM_2_59_port, IN4 => n2636, Q => n3065);
   U3082 : AO22X2 port map( IN1 => RAM_3_7_port, IN2 => n2549, IN3 => 
                           RAM_2_7_port, IN4 => n2624, Q => n2857);
   U3083 : AO22X2 port map( IN1 => RAM_11_1_port, IN2 => n3453, IN3 => 
                           RAM_10_1_port, IN4 => n2655, Q => n2831);
   U3084 : AO22X2 port map( IN1 => RAM_11_100_port, IN2 => n3454, IN3 => n2657,
                           IN4 => RAM_10_100_port, Q => n3227);
   U3085 : AO22X2 port map( IN1 => RAM_11_77_port, IN2 => n3455, IN3 => n2661, 
                           IN4 => RAM_10_77_port, Q => n3135);
   U3086 : AO22X2 port map( IN1 => RAM_11_114_port, IN2 => n2501, IN3 => 
                           RAM_10_114_port, IN4 => n2661, Q => n3287);
   U3087 : AO22X2 port map( IN1 => RAM_11_2_port, IN2 => n2501, IN3 => 
                           RAM_10_2_port, IN4 => n2659, Q => n2835);
   U3088 : AO22X2 port map( IN1 => n3453, IN2 => RAM_11_59_port, IN3 => 
                           RAM_10_59_port, IN4 => n2660, Q => n3063);
   U3089 : AO22X2 port map( IN1 => n3460, IN2 => RAM_11_25_port, IN3 => n2651, 
                           IN4 => RAM_10_25_port, Q => n2927);
   U3090 : OR4X2 port map( IN1 => n4184, IN2 => n4183, IN3 => n4182, IN4 => 
                           n4181, Q => RAMDOUT2(88));
   U3091 : AND2X4 port map( IN1 => n2797, IN2 => n2202, Q => n2742);
   U3092 : AND2X4 port map( IN1 => n2797, IN2 => n2202, Q => n2743);
   U3093 : AND2X4 port map( IN1 => n2797, IN2 => n2202, Q => n3353);
   U3094 : NAND4X0 port map( IN1 => n2744, IN2 => n2745, IN3 => n2746, IN4 => 
                           n2747, QN => RAMDOUT1(120));
   U3095 : AOI221X1 port map( IN1 => RAM_8_120_port, IN2 => n3419, IN3 => 
                           RAM_9_120_port, IN4 => n3360, IN5 => n3311, QN => 
                           n2744);
   U3096 : AOI221X1 port map( IN1 => RAM_12_120_port, IN2 => n2449, IN3 => 
                           RAM_13_120_port, IN4 => n3373, IN5 => n3312, QN => 
                           n2745);
   U3097 : AOI221X1 port map( IN1 => RAM_0_120_port, IN2 => n2167, IN3 => 
                           RAM_1_120_port, IN4 => n2157, IN5 => n3313, QN => 
                           n2746);
   U3098 : AOI221X1 port map( IN1 => RAM_4_120_port, IN2 => n3406, IN3 => 
                           RAM_5_120_port, IN4 => n2495, IN5 => n3314, QN => 
                           n2747);
   U3099 : AO22X2 port map( IN1 => RAM_7_98_port, IN2 => n2525, IN3 => 
                           RAM_6_98_port, IN4 => n2135, Q => n3222);
   U3100 : AO22X2 port map( IN1 => RAM_7_45_port, IN2 => n2517, IN3 => 
                           RAM_6_45_port, IN4 => n2150, Q => n3010);
   U3101 : AO22X2 port map( IN1 => RAM_7_64_port, IN2 => n2525, IN3 => 
                           RAM_6_64_port, IN4 => n2135, Q => n3086);
   U3102 : AO22X2 port map( IN1 => RAM_7_75_port, IN2 => n2524, IN3 => 
                           RAM_6_75_port, IN4 => n2148, Q => n3130);
   U3103 : AO22X2 port map( IN1 => RAM_7_38_port, IN2 => n2528, IN3 => 
                           RAM_6_38_port, IN4 => n2137, Q => n2982);
   U3104 : AO22X2 port map( IN1 => RAM_7_59_port, IN2 => n2394, IN3 => 
                           RAM_6_59_port, IN4 => n2142, Q => n3066);
   U3105 : AO22X2 port map( IN1 => RAM_7_127_port, IN2 => n2528, IN3 => 
                           RAM_6_127_port, IN4 => n2134, Q => n3355);
   U3106 : AO22X2 port map( IN1 => RAM_7_70_port, IN2 => n2522, IN3 => 
                           RAM_6_70_port, IN4 => n2138, Q => n3110);
   U3107 : AO22X2 port map( IN1 => RAM_7_51_port, IN2 => n2520, IN3 => 
                           RAM_6_51_port, IN4 => n2141, Q => n3034);
   U3108 : AO22X2 port map( IN1 => RAM_7_81_port, IN2 => n2519, IN3 => 
                           RAM_6_81_port, IN4 => n2150, Q => n3154);
   U3109 : AO22X2 port map( IN1 => RAM_7_73_port, IN2 => n2524, IN3 => 
                           RAM_6_73_port, IN4 => n2136, Q => n3122);
   U3110 : AO22X2 port map( IN1 => RAM_7_23_port, IN2 => n2521, IN3 => 
                           RAM_6_23_port, IN4 => n2140, Q => n2922);
   U3111 : AO22X2 port map( IN1 => RAM_7_115_port, IN2 => n2530, IN3 => 
                           RAM_6_115_port, IN4 => n2143, Q => n3294);
   U3112 : AO22X2 port map( IN1 => RAM_7_29_port, IN2 => n2520, IN3 => 
                           RAM_6_29_port, IN4 => n2138, Q => n2946);
   U3113 : AO22X2 port map( IN1 => RAM_7_39_port, IN2 => n2516, IN3 => 
                           RAM_6_39_port, IN4 => n2146, Q => n2986);
   U3114 : AO22X2 port map( IN1 => RAM_7_63_port, IN2 => n2513, IN3 => 
                           RAM_6_63_port, IN4 => n2144, Q => n3082);
   U3115 : AO22X2 port map( IN1 => RAM_7_52_port, IN2 => n2530, IN3 => 
                           RAM_6_52_port, IN4 => n2141, Q => n3038);
   U3116 : AO22X2 port map( IN1 => RAM_7_11_port, IN2 => n2522, IN3 => 
                           RAM_6_11_port, IN4 => n2147, Q => n2874);
   U3117 : AO22X2 port map( IN1 => RAM_7_111_port, IN2 => n2521, IN3 => 
                           RAM_6_111_port, IN4 => n2148, Q => n3274);
   U3118 : AO22X2 port map( IN1 => RAM_7_22_port, IN2 => n2514, IN3 => 
                           RAM_6_22_port, IN4 => n2142, Q => n2918);
   U3119 : AND2X4 port map( IN1 => n2797, IN2 => n2821, Q => n2748);
   U3120 : AND2X4 port map( IN1 => n2797, IN2 => n2821, Q => n3343);
   U3121 : OR4X2 port map( IN1 => n4464, IN2 => n4463, IN3 => n4462, IN4 => 
                           n4461, Q => RAMDOUT2(123));
   U3122 : NAND4X0 port map( IN1 => n2749, IN2 => n2750, IN3 => n2751, IN4 => 
                           n2752, QN => RAMDOUT1(27));
   U3123 : AOI221X2 port map( IN1 => RAM_8_27_port, IN2 => n3419, IN3 => 
                           RAM_9_27_port, IN4 => n3369, IN5 => n2935, QN => 
                           n2749);
   U3124 : AOI221X1 port map( IN1 => RAM_12_27_port, IN2 => n2449, IN3 => 
                           RAM_13_27_port, IN4 => n3378, IN5 => n2936, QN => 
                           n2750);
   U3125 : AOI221X1 port map( IN1 => RAM_0_27_port, IN2 => n2162, IN3 => 
                           RAM_1_27_port, IN4 => n3383, IN5 => n2937, QN => 
                           n2751);
   U3126 : AOI221X2 port map( IN1 => RAM_4_27_port, IN2 => n3406, IN3 => 
                           RAM_5_27_port, IN4 => n3397, IN5 => n2938, QN => 
                           n2752);
   U3127 : NAND4X0 port map( IN1 => n2755, IN2 => n2753, IN3 => n2754, IN4 => 
                           n2756, QN => RAMDOUT1(81));
   U3128 : AOI221X1 port map( IN1 => RAM_8_81_port, IN2 => n3420, IN3 => 
                           RAM_9_81_port, IN4 => n3363, IN5 => n3151, QN => 
                           n2753);
   U3129 : AOI221X1 port map( IN1 => RAM_12_81_port, IN2 => n2458, IN3 => 
                           RAM_13_81_port, IN4 => n3371, IN5 => n3152, QN => 
                           n2754);
   U3130 : AOI221X1 port map( IN1 => RAM_0_81_port, IN2 => n2162, IN3 => 
                           RAM_1_81_port, IN4 => n2121, IN5 => n3153, QN => 
                           n2755);
   U3131 : AOI221X2 port map( IN1 => RAM_4_81_port, IN2 => n3408, IN3 => 
                           RAM_5_81_port, IN4 => n2494, IN5 => n3154, QN => 
                           n2756);
   U3132 : AO22X2 port map( IN1 => RAM_15_105_port, IN2 => n3441, IN3 => 
                           RAM_14_105_port, IN4 => n2330, Q => n3248);
   U3133 : AO22X2 port map( IN1 => RAM_15_8_port, IN2 => n3439, IN3 => 
                           RAM_14_8_port, IN4 => n2335, Q => n2860);
   U3134 : AO22X2 port map( IN1 => RAM_15_6_port, IN2 => n3436, IN3 => 
                           RAM_14_6_port, IN4 => n2321, Q => n2852);
   U3135 : AO22X2 port map( IN1 => RAM_15_111_port, IN2 => n3439, IN3 => 
                           RAM_14_111_port, IN4 => n2321, Q => n3272);
   U3136 : AO22X2 port map( IN1 => RAM_15_84_port, IN2 => n3436, IN3 => 
                           RAM_14_84_port, IN4 => n2323, Q => n3164);
   U3137 : AO22X2 port map( IN1 => RAM_15_22_port, IN2 => n3446, IN3 => 
                           RAM_14_22_port, IN4 => n2333, Q => n2916);
   U3138 : AO22X2 port map( IN1 => RAM_15_13_port, IN2 => n3444, IN3 => 
                           RAM_14_13_port, IN4 => n2330, Q => n2880);
   U3139 : AO22X2 port map( IN1 => RAM_15_63_port, IN2 => n3434, IN3 => 
                           RAM_14_63_port, IN4 => n2339, Q => n3080);
   U3140 : AO22X2 port map( IN1 => RAM_15_37_port, IN2 => n3440, IN3 => 
                           RAM_14_37_port, IN4 => n2325, Q => n2976);
   U3141 : AO22X2 port map( IN1 => RAM_15_20_port, IN2 => n3435, IN3 => 
                           RAM_14_20_port, IN4 => n2321, Q => n2908);
   U3142 : AO22X2 port map( IN1 => RAM_15_106_port, IN2 => n3436, IN3 => 
                           RAM_14_106_port, IN4 => n2338, Q => n3252);
   U3143 : AO22X2 port map( IN1 => RAM_15_3_port, IN2 => n3439, IN3 => 
                           RAM_14_3_port, IN4 => n2329, Q => n2840);
   U3144 : AO22X2 port map( IN1 => RAM_15_117_port, IN2 => n3432, IN3 => 
                           RAM_14_117_port, IN4 => n2324, Q => n3300);
   U3145 : AO22X2 port map( IN1 => RAM_15_123_port, IN2 => n3440, IN3 => 
                           RAM_14_123_port, IN4 => n2321, Q => n3324);
   U3146 : AO22X2 port map( IN1 => RAM_15_122_port, IN2 => n3440, IN3 => 
                           RAM_14_122_port, IN4 => n2326, Q => n3320);
   U3147 : AO22X2 port map( IN1 => RAM_15_95_port, IN2 => n3441, IN3 => 
                           RAM_14_95_port, IN4 => n2325, Q => n3208);
   U3148 : NAND4X0 port map( IN1 => n2757, IN2 => n2758, IN3 => n2759, IN4 => 
                           n2760, QN => RAMDOUT1(26));
   U3149 : AOI221X1 port map( IN1 => RAM_8_26_port, IN2 => n3416, IN3 => 
                           RAM_9_26_port, IN4 => n3364, IN5 => n2931, QN => 
                           n2757);
   U3150 : AOI221X1 port map( IN1 => RAM_4_26_port, IN2 => n3404, IN3 => 
                           RAM_5_26_port, IN4 => n3391, IN5 => n2934, QN => 
                           n2760);
   U3151 : AO22X2 port map( IN1 => RAM_3_45_port, IN2 => n2552, IN3 => 
                           RAM_2_45_port, IN4 => n2640, Q => n3009);
   U3152 : AO22X2 port map( IN1 => RAM_3_48_port, IN2 => n2479, IN3 => 
                           RAM_2_48_port, IN4 => n2632, Q => n3021);
   U3153 : AO22X2 port map( IN1 => RAM_3_53_port, IN2 => n2546, IN3 => 
                           RAM_2_53_port, IN4 => n2624, Q => n3041);
   U3154 : AO22X2 port map( IN1 => RAM_3_18_port, IN2 => n2546, IN3 => 
                           RAM_2_18_port, IN4 => n2099, Q => n2901);
   U3155 : AO22X2 port map( IN1 => RAM_3_102_port, IN2 => n2479, IN3 => 
                           RAM_2_102_port, IN4 => n2111, Q => n3237);
   U3156 : AO22X2 port map( IN1 => RAM_3_83_port, IN2 => n2538, IN3 => 
                           RAM_2_83_port, IN4 => n2099, Q => n3161);
   U3157 : AO22X2 port map( IN1 => RAM_3_76_port, IN2 => n2544, IN3 => n2638, 
                           IN4 => RAM_2_76_port, Q => n3133);
   U3158 : AO22X2 port map( IN1 => RAM_3_90_port, IN2 => n2399, IN3 => 
                           RAM_2_90_port, IN4 => n2641, Q => n3189);
   U3159 : AO22X2 port map( IN1 => RAM_3_66_port, IN2 => n2539, IN3 => n2644, 
                           IN4 => RAM_2_66_port, Q => n3093);
   U3160 : AO22X2 port map( IN1 => RAM_3_85_port, IN2 => n2545, IN3 => 
                           RAM_2_85_port, IN4 => n2631, Q => n3169);
   U3161 : AO22X2 port map( IN1 => RAM_3_27_port, IN2 => n2399, IN3 => 
                           RAM_2_27_port, IN4 => n2626, Q => n2937);
   U3162 : AO22X2 port map( IN1 => RAM_3_88_port, IN2 => n2470, IN3 => 
                           RAM_2_88_port, IN4 => n2623, Q => n3181);
   U3163 : AO22X2 port map( IN1 => RAM_3_40_port, IN2 => n2538, IN3 => 
                           RAM_2_40_port, IN4 => n2630, Q => n2989);
   U3164 : AO22X2 port map( IN1 => RAM_3_113_port, IN2 => n2553, IN3 => 
                           RAM_2_113_port, IN4 => n2627, Q => n3285);
   U3165 : AO22X2 port map( IN1 => RAM_3_24_port, IN2 => n2550, IN3 => 
                           RAM_2_24_port, IN4 => n2638, Q => n2925);
   U3166 : AO22X2 port map( IN1 => RAM_3_14_port, IN2 => n2541, IN3 => 
                           RAM_2_14_port, IN4 => n2623, Q => n2885);
   U3167 : AO22X2 port map( IN1 => RAM_3_23_port, IN2 => n2540, IN3 => 
                           RAM_2_23_port, IN4 => n2111, Q => n2921);
   U3168 : AO22X2 port map( IN1 => RAM_3_123_port, IN2 => n2542, IN3 => 
                           RAM_2_123_port, IN4 => n2635, Q => n3325);
   U3169 : AO22X2 port map( IN1 => RAM_3_93_port, IN2 => n2544, IN3 => n2631, 
                           IN4 => RAM_2_93_port, Q => n3201);
   U3170 : AO22X2 port map( IN1 => RAM_3_101_port, IN2 => n2541, IN3 => 
                           RAM_2_101_port, IN4 => n2639, Q => n3233);
   U3171 : AO22X2 port map( IN1 => RAM_3_92_port, IN2 => n2551, IN3 => n2631, 
                           IN4 => RAM_2_92_port, Q => n3197);
   U3172 : AO22X2 port map( IN1 => RAM_3_25_port, IN2 => n2539, IN3 => 
                           RAM_2_25_port, IN4 => n2632, Q => n2929);
   U3173 : NAND4X0 port map( IN1 => n2761, IN2 => n2762, IN3 => n2763, IN4 => 
                           n2764, QN => RAMDOUT1(2));
   U3174 : AOI221X1 port map( IN1 => RAM_8_2_port, IN2 => n3421, IN3 => 
                           RAM_9_2_port, IN4 => n2493, IN5 => n2835, QN => 
                           n2761);
   U3175 : AOI221X1 port map( IN1 => RAM_12_2_port, IN2 => n2446, IN3 => 
                           RAM_13_2_port, IN4 => n2489, IN5 => n2836, QN => 
                           n2762);
   U3176 : AOI221X1 port map( IN1 => RAM_0_2_port, IN2 => n2173, IN3 => 
                           RAM_1_2_port, IN4 => n3390, IN5 => n2837, QN => 
                           n2763);
   U3177 : AOI221X1 port map( IN1 => RAM_4_2_port, IN2 => n3402, IN3 => 
                           RAM_5_2_port, IN4 => n3394, IN5 => n2838, QN => 
                           n2764);
   U3178 : AO22X2 port map( IN1 => RAM_15_88_port, IN2 => n3438, IN3 => 
                           RAM_14_88_port, IN4 => n2326, Q => n3180);
   U3179 : AO22X2 port map( IN1 => RAM_15_32_port, IN2 => n3440, IN3 => 
                           RAM_14_32_port, IN4 => n2332, Q => n2956);
   U3180 : AO22X2 port map( IN1 => RAM_15_42_port, IN2 => n3435, IN3 => 
                           RAM_14_42_port, IN4 => n2336, Q => n2996);
   U3181 : AO22X2 port map( IN1 => RAM_15_55_port, IN2 => n3445, IN3 => 
                           RAM_14_55_port, IN4 => n2323, Q => n3048);
   U3182 : AO22X2 port map( IN1 => RAM_15_12_port, IN2 => n3445, IN3 => 
                           RAM_14_12_port, IN4 => n2322, Q => n2876);
   U3183 : AO22X2 port map( IN1 => RAM_15_16_port, IN2 => n3433, IN3 => 
                           RAM_14_16_port, IN4 => n2337, Q => n2892);
   U3184 : AO22X2 port map( IN1 => RAM_15_72_port, IN2 => n3439, IN3 => 
                           RAM_14_72_port, IN4 => n2328, Q => n3116);
   U3185 : AO22X2 port map( IN1 => RAM_15_116_port, IN2 => n3438, IN3 => 
                           RAM_14_116_port, IN4 => n2337, Q => n3296);
   U3186 : AO22X2 port map( IN1 => RAM_15_67_port, IN2 => n3440, IN3 => 
                           RAM_14_67_port, IN4 => n2338, Q => n3096);
   U3187 : AO22X2 port map( IN1 => RAM_15_25_port, IN2 => n3432, IN3 => 
                           RAM_14_25_port, IN4 => n2322, Q => n2928);
   U3188 : AO22X2 port map( IN1 => RAM_15_90_port, IN2 => n3434, IN3 => 
                           RAM_14_90_port, IN4 => n2320, Q => n3188);
   U3189 : AO22X2 port map( IN1 => RAM_15_54_port, IN2 => n3432, IN3 => 
                           RAM_14_54_port, IN4 => n2325, Q => n3044);
   U3190 : AO22X2 port map( IN1 => RAM_15_62_port, IN2 => n3437, IN3 => 
                           RAM_14_62_port, IN4 => n2328, Q => n3076);
   U3191 : AO22X2 port map( IN1 => RAM_15_64_port, IN2 => n3436, IN3 => 
                           RAM_14_64_port, IN4 => n2337, Q => n3084);
   U3192 : AO22X2 port map( IN1 => RAM_15_15_port, IN2 => n3438, IN3 => 
                           RAM_14_15_port, IN4 => n2329, Q => n2888);
   U3193 : AO22X2 port map( IN1 => RAM_15_83_port, IN2 => n3445, IN3 => 
                           RAM_14_83_port, IN4 => n2328, Q => n3160);
   U3194 : AO22X2 port map( IN1 => RAM_15_115_port, IN2 => n3446, IN3 => 
                           RAM_14_115_port, IN4 => n2327, Q => n3292);
   U3195 : AO22X2 port map( IN1 => RAM_15_75_port, IN2 => n3446, IN3 => 
                           RAM_14_75_port, IN4 => n2327, Q => n3128);
   U3196 : AO22X2 port map( IN1 => RAM_15_107_port, IN2 => n3441, IN3 => 
                           RAM_14_107_port, IN4 => n2320, Q => n3256);
   U3197 : AO22X2 port map( IN1 => RAM_15_80_port, IN2 => n3437, IN3 => 
                           RAM_14_80_port, IN4 => n2329, Q => n3148);
   U3198 : AO22X2 port map( IN1 => RAM_15_69_port, IN2 => n3438, IN3 => 
                           RAM_14_69_port, IN4 => n2330, Q => n3104);
   U3199 : AO22X2 port map( IN1 => RAM_15_31_port, IN2 => n3444, IN3 => 
                           RAM_14_31_port, IN4 => n2330, Q => n2952);
   U3200 : NAND4X0 port map( IN1 => n2765, IN2 => n2766, IN3 => n2767, IN4 => 
                           n2768, QN => RAMDOUT1(123));
   U3201 : AOI221X1 port map( IN1 => RAM_8_123_port, IN2 => n3423, IN3 => 
                           RAM_9_123_port, IN4 => n3364, IN5 => n3323, QN => 
                           n2765);
   U3202 : AOI221X1 port map( IN1 => RAM_12_123_port, IN2 => n2459, IN3 => 
                           RAM_13_123_port, IN4 => n3375, IN5 => n3324, QN => 
                           n2766);
   U3203 : AOI221X1 port map( IN1 => RAM_0_123_port, IN2 => n2159, IN3 => 
                           RAM_1_123_port, IN4 => n3383, IN5 => n3325, QN => 
                           n2767);
   U3204 : AOI221X1 port map( IN1 => RAM_4_123_port, IN2 => n3448, IN3 => 
                           RAM_5_123_port, IN4 => n3399, IN5 => n3326, QN => 
                           n2768);
   U3205 : AOI221X1 port map( IN1 => RAM_8_92_port, IN2 => n3416, IN3 => 
                           RAM_9_92_port, IN4 => n3360, IN5 => n3195, QN => 
                           n2781);
   U3206 : AOI221X1 port map( IN1 => RAM_8_68_port, IN2 => n3425, IN3 => 
                           RAM_9_68_port, IN4 => n3363, IN5 => n3099, QN => 
                           n2785);
   U3207 : AO22X2 port map( IN1 => RAM_15_39_port, IN2 => n3434, IN3 => 
                           RAM_14_39_port, IN4 => n2333, Q => n2984);
   U3208 : AO22X2 port map( IN1 => RAM_15_36_port, IN2 => n3445, IN3 => 
                           RAM_14_36_port, IN4 => n2331, Q => n2972);
   U3209 : AO22X2 port map( IN1 => RAM_15_23_port, IN2 => n3433, IN3 => 
                           RAM_14_23_port, IN4 => n2338, Q => n2920);
   U3210 : AO22X2 port map( IN1 => RAM_15_21_port, IN2 => n3434, IN3 => 
                           RAM_14_21_port, IN4 => n2330, Q => n2912);
   U3211 : AO22X2 port map( IN1 => RAM_15_79_port, IN2 => n3432, IN3 => 
                           RAM_14_79_port, IN4 => n2332, Q => n3144);
   U3212 : AO22X2 port map( IN1 => RAM_15_100_port, IN2 => n3441, IN3 => 
                           RAM_14_100_port, IN4 => n2336, Q => n3228);
   U3213 : AO22X2 port map( IN1 => RAM_15_85_port, IN2 => n3433, IN3 => 
                           RAM_14_85_port, IN4 => n2327, Q => n3168);
   U3214 : AO22X2 port map( IN1 => RAM_15_29_port, IN2 => n3444, IN3 => 
                           RAM_14_29_port, IN4 => n2320, Q => n2944);
   U3215 : AO22X2 port map( IN1 => RAM_15_1_port, IN2 => n3441, IN3 => 
                           RAM_14_1_port, IN4 => n2336, Q => n2832);
   U3216 : AO22X2 port map( IN1 => RAM_15_46_port, IN2 => n3437, IN3 => 
                           RAM_14_46_port, IN4 => n2339, Q => n3012);
   U3217 : AO22X2 port map( IN1 => RAM_15_73_port, IN2 => n3444, IN3 => 
                           RAM_14_73_port, IN4 => n2333, Q => n3120);
   U3218 : AO22X2 port map( IN1 => RAM_15_10_port, IN2 => n3435, IN3 => 
                           RAM_14_10_port, IN4 => n2334, Q => n2868);
   U3219 : AO22X2 port map( IN1 => RAM_15_52_port, IN2 => n3437, IN3 => 
                           RAM_14_52_port, IN4 => n2324, Q => n3036);
   U3220 : AO22X2 port map( IN1 => RAM_15_17_port, IN2 => n3441, IN3 => 
                           RAM_14_17_port, IN4 => n2322, Q => n2896);
   U3221 : AO22X2 port map( IN1 => RAM_15_114_port, IN2 => n3435, IN3 => 
                           RAM_14_114_port, IN4 => n2335, Q => n3288);
   U3222 : AO22X2 port map( IN1 => RAM_15_74_port, IN2 => n3432, IN3 => 
                           RAM_14_74_port, IN4 => n2329, Q => n3124);
   U3223 : AO22X2 port map( IN1 => RAM_15_125_port, IN2 => n3440, IN3 => 
                           RAM_14_125_port, IN4 => n2323, Q => n3332);
   U3224 : AO22X2 port map( IN1 => RAM_15_26_port, IN2 => n3434, IN3 => 
                           RAM_14_26_port, IN4 => n2324, Q => n2932);
   U3225 : AO22X2 port map( IN1 => RAM_15_33_port, IN2 => n3439, IN3 => 
                           RAM_14_33_port, IN4 => n2328, Q => n2960);
   U3226 : AO22X2 port map( IN1 => RAM_15_43_port, IN2 => n3435, IN3 => 
                           RAM_14_43_port, IN4 => n2333, Q => n3000);
   U3227 : AO22X2 port map( IN1 => RAM_15_48_port, IN2 => n3445, IN3 => 
                           RAM_14_48_port, IN4 => n2325, Q => n3020);
   U3228 : AO22X2 port map( IN1 => RAM_15_9_port, IN2 => n3446, IN3 => 
                           RAM_14_9_port, IN4 => n2332, Q => n2864);
   U3229 : AO22X2 port map( IN1 => RAM_15_124_port, IN2 => n3438, IN3 => 
                           RAM_14_124_port, IN4 => n2333, Q => n3328);
   U3230 : AO22X2 port map( IN1 => RAM_15_93_port, IN2 => n3435, IN3 => 
                           RAM_14_93_port, IN4 => n2325, Q => n3200);
   U3231 : AO22X2 port map( IN1 => RAM_15_121_port, IN2 => n3432, IN3 => 
                           RAM_14_121_port, IN4 => n2325, Q => n3316);
   U3232 : AO22X2 port map( IN1 => RAM_15_126_port, IN2 => n3436, IN3 => 
                           RAM_14_126_port, IN4 => n2331, Q => n3336);
   U3233 : AO22X2 port map( IN1 => RAM_15_2_port, IN2 => n3434, IN3 => 
                           RAM_14_2_port, IN4 => n2327, Q => n2836);
   U3234 : AO22X2 port map( IN1 => RAM_11_54_port, IN2 => n3449, IN3 => 
                           RAM_10_54_port, IN4 => n2666, Q => n3043);
   U3235 : AO22X2 port map( IN1 => RAM_11_12_port, IN2 => n3455, IN3 => 
                           RAM_10_12_port, IN4 => n2653, Q => n2875);
   U3236 : AO22X2 port map( IN1 => RAM_11_23_port, IN2 => n3453, IN3 => 
                           RAM_10_23_port, IN4 => n2663, Q => n2919);
   U3237 : AO22X2 port map( IN1 => RAM_11_20_port, IN2 => n3450, IN3 => n2650, 
                           IN4 => RAM_10_20_port, Q => n2907);
   U3238 : AO22X2 port map( IN1 => RAM_11_69_port, IN2 => n3459, IN3 => n2480, 
                           IN4 => RAM_10_69_port, Q => n3103);
   U3239 : AO22X2 port map( IN1 => RAM_11_88_port, IN2 => n3457, IN3 => 
                           RAM_10_88_port, IN4 => n2664, Q => n3179);
   U3240 : AO22X2 port map( IN1 => RAM_11_53_port, IN2 => n2504, IN3 => n2480, 
                           IN4 => RAM_10_53_port, Q => n3039);
   U3241 : AO22X2 port map( IN1 => RAM_11_18_port, IN2 => n3449, IN3 => n2373, 
                           IN4 => RAM_10_18_port, Q => n2899);
   U3242 : AO22X2 port map( IN1 => RAM_11_4_port, IN2 => n2231, IN3 => n2373, 
                           IN4 => RAM_10_4_port, Q => n2843);
   U3243 : AO22X2 port map( IN1 => RAM_11_80_port, IN2 => n3449, IN3 => 
                           RAM_10_80_port, IN4 => n2654, Q => n3147);
   U3244 : AO22X2 port map( IN1 => RAM_11_26_port, IN2 => n3454, IN3 => n2654, 
                           IN4 => RAM_10_26_port, Q => n2931);
   U3245 : AO22X2 port map( IN1 => RAM_11_126_port, IN2 => n3462, IN3 => n2654,
                           IN4 => RAM_10_126_port, Q => n3335);
   U3246 : AO22X2 port map( IN1 => RAM_11_29_port, IN2 => n3458, IN3 => n2665, 
                           IN4 => RAM_10_29_port, Q => n2943);
   U3247 : AO22X2 port map( IN1 => RAM_11_118_port, IN2 => n3453, IN3 => 
                           RAM_10_118_port, IN4 => n2657, Q => n3303);
   U3248 : AO22X2 port map( IN1 => RAM_11_61_port, IN2 => n3461, IN3 => 
                           RAM_10_61_port, IN4 => n2461, Q => n3071);
   U3249 : AO22X2 port map( IN1 => RAM_11_76_port, IN2 => n3453, IN3 => 
                           RAM_10_76_port, IN4 => n2667, Q => n3131);
   U3250 : AO22X2 port map( IN1 => RAM_11_119_port, IN2 => n3458, IN3 => 
                           RAM_10_119_port, IN4 => n2653, Q => n3307);
   U3251 : AO22X2 port map( IN1 => RAM_11_124_port, IN2 => n3454, IN3 => 
                           RAM_10_124_port, IN4 => n2660, Q => n3327);
   U3252 : AO22X2 port map( IN1 => RAM_11_84_port, IN2 => n2501, IN3 => 
                           RAM_10_84_port, IN4 => n2651, Q => n3163);
   U3253 : AO22X2 port map( IN1 => RAM_11_120_port, IN2 => n3452, IN3 => 
                           RAM_10_120_port, IN4 => n2191, Q => n3311);
   U3254 : AO22X2 port map( IN1 => RAM_11_22_port, IN2 => n2504, IN3 => 
                           RAM_10_22_port, IN4 => n2467, Q => n2915);
   U3255 : AO22X2 port map( IN1 => RAM_3_20_port, IN2 => n2469, IN3 => n7, IN4 
                           => RAM_2_20_port, Q => n2909);
   U3256 : NAND4X0 port map( IN1 => n2769, IN2 => n2771, IN3 => n2770, IN4 => 
                           n2772, QN => RAMDOUT1(93));
   U3257 : AOI221X1 port map( IN1 => RAM_8_93_port, IN2 => n3420, IN3 => 
                           RAM_9_93_port, IN4 => n3362, IN5 => n3199, QN => 
                           n2769);
   U3258 : AOI221X1 port map( IN1 => RAM_12_93_port, IN2 => n2460, IN3 => 
                           RAM_13_93_port, IN4 => n2489, IN5 => n3200, QN => 
                           n2770);
   U3259 : AOI221X1 port map( IN1 => RAM_0_93_port, IN2 => n2161, IN3 => 
                           RAM_1_93_port, IN4 => n3387, IN5 => n3201, QN => 
                           n2771);
   U3260 : AOI221X2 port map( IN1 => RAM_4_93_port, IN2 => n3407, IN3 => 
                           RAM_5_93_port, IN4 => n3397, IN5 => n3202, QN => 
                           n2772);
   U3261 : NAND4X0 port map( IN1 => n2773, IN2 => n2774, IN3 => n2775, IN4 => 
                           n2776, QN => RAMDOUT1(108));
   U3262 : AOI221X1 port map( IN1 => RAM_8_108_port, IN2 => n3424, IN3 => 
                           RAM_9_108_port, IN4 => n3364, IN5 => n3259, QN => 
                           n2773);
   U3263 : AOI221X1 port map( IN1 => RAM_12_108_port, IN2 => n2445, IN3 => 
                           RAM_13_108_port, IN4 => n3371, IN5 => n3260, QN => 
                           n2774);
   U3264 : AOI221X1 port map( IN1 => RAM_0_108_port, IN2 => n2169, IN3 => 
                           RAM_1_108_port, IN4 => n2491, IN5 => n3261, QN => 
                           n2775);
   U3265 : AOI221X1 port map( IN1 => RAM_4_108_port, IN2 => n3410, IN3 => 
                           RAM_5_108_port, IN4 => n3396, IN5 => n3262, QN => 
                           n2776);
   U3266 : AO22X2 port map( IN1 => RAM_15_120_port, IN2 => n3445, IN3 => 
                           RAM_14_120_port, IN4 => n2339, Q => n3312);
   U3267 : NAND4X0 port map( IN1 => n2777, IN2 => n2778, IN3 => n2779, IN4 => 
                           n2780, QN => RAMDOUT1(67));
   U3268 : AOI221X1 port map( IN1 => RAM_8_67_port, IN2 => n3422, IN3 => 
                           RAM_9_67_port, IN4 => n2493, IN5 => n3095, QN => 
                           n2777);
   U3269 : AOI221X1 port map( IN1 => RAM_12_67_port, IN2 => n2452, IN3 => 
                           RAM_13_67_port, IN4 => n3373, IN5 => n3096, QN => 
                           n2778);
   U3270 : AOI221X1 port map( IN1 => RAM_0_67_port, IN2 => n2169, IN3 => 
                           RAM_1_67_port, IN4 => n3387, IN5 => n3097, QN => 
                           n2779);
   U3271 : AOI221X1 port map( IN1 => RAM_4_67_port, IN2 => n3448, IN3 => 
                           RAM_5_67_port, IN4 => n3393, IN5 => n3098, QN => 
                           n2780);
   U3272 : NAND4X0 port map( IN1 => n2781, IN2 => n2782, IN3 => n2783, IN4 => 
                           n2784, QN => RAMDOUT1(92));
   U3273 : AOI221X1 port map( IN1 => RAM_12_92_port, IN2 => n2460, IN3 => 
                           RAM_13_92_port, IN4 => n3372, IN5 => n3196, QN => 
                           n2782);
   U3274 : AOI221X1 port map( IN1 => RAM_0_92_port, IN2 => n2165, IN3 => 
                           RAM_1_92_port, IN4 => n3387, IN5 => n3197, QN => 
                           n2783);
   U3275 : AOI221X2 port map( IN1 => RAM_4_92_port, IN2 => n3408, IN3 => 
                           RAM_5_92_port, IN4 => n3397, IN5 => n3198, QN => 
                           n2784);
   U3276 : NAND4X0 port map( IN1 => n2785, IN2 => n2786, IN3 => n2787, IN4 => 
                           n2788, QN => RAMDOUT1(68));
   U3277 : AOI221X1 port map( IN1 => RAM_12_68_port, IN2 => n2460, IN3 => 
                           RAM_13_68_port, IN4 => n3377, IN5 => n3100, QN => 
                           n2786);
   U3278 : AOI221X2 port map( IN1 => RAM_4_68_port, IN2 => n3409, IN3 => 
                           RAM_5_68_port, IN4 => n3399, IN5 => n3102, QN => 
                           n2788);
   U3279 : NAND4X0 port map( IN1 => n2789, IN2 => n2790, IN3 => n2791, IN4 => 
                           n2792, QN => RAMDOUT1(6));
   U3280 : AOI221X1 port map( IN1 => RAM_8_6_port, IN2 => n3423, IN3 => 
                           RAM_9_6_port, IN4 => n2493, IN5 => n2851, QN => 
                           n2789);
   U3281 : AOI221X1 port map( IN1 => RAM_12_6_port, IN2 => n2453, IN3 => 
                           RAM_13_6_port, IN4 => n3376, IN5 => n2852, QN => 
                           n2790);
   U3282 : AOI221X1 port map( IN1 => RAM_0_6_port, IN2 => n2160, IN3 => 
                           RAM_1_6_port, IN4 => n3390, IN5 => n2853, QN => 
                           n2791);
   U3283 : AOI221X1 port map( IN1 => RAM_4_6_port, IN2 => n3406, IN3 => 
                           RAM_5_6_port, IN4 => n3391, IN5 => n2854, QN => 
                           n2792);
   U3284 : NAND4X0 port map( IN1 => n2793, IN2 => n2794, IN3 => n2795, IN4 => 
                           n2796, QN => RAMDOUT1(98));
   U3285 : AOI221X1 port map( IN1 => RAM_8_98_port, IN2 => n3425, IN3 => 
                           RAM_9_98_port, IN4 => n3368, IN5 => n3219, QN => 
                           n2793);
   U3286 : AOI221X1 port map( IN1 => RAM_12_98_port, IN2 => n2452, IN3 => 
                           RAM_13_98_port, IN4 => n3372, IN5 => n3220, QN => 
                           n2794);
   U3287 : AOI221X1 port map( IN1 => RAM_0_98_port, IN2 => n2161, IN3 => 
                           RAM_1_98_port, IN4 => n3384, IN5 => n3221, QN => 
                           n2795);
   U3288 : AOI221X2 port map( IN1 => RAM_4_98_port, IN2 => n3409, IN3 => 
                           RAM_5_98_port, IN4 => n3400, IN5 => n3222, QN => 
                           n2796);
   U3289 : NAND4X0 port map( IN1 => n2798, IN2 => n2799, IN3 => n2800, IN4 => 
                           n2801, QN => RAMDOUT1(121));
   U3290 : AOI221X1 port map( IN1 => RAM_8_121_port, IN2 => n3424, IN3 => 
                           RAM_9_121_port, IN4 => n3367, IN5 => n3315, QN => 
                           n2798);
   U3291 : AOI221X1 port map( IN1 => RAM_12_121_port, IN2 => n2447, IN3 => 
                           RAM_13_121_port, IN4 => n3374, IN5 => n3316, QN => 
                           n2799);
   U3292 : AOI221X1 port map( IN1 => RAM_0_121_port, IN2 => n2164, IN3 => 
                           RAM_1_121_port, IN4 => n3389, IN5 => n3317, QN => 
                           n2800);
   U3293 : NAND4X0 port map( IN1 => n2802, IN2 => n2803, IN3 => n2804, IN4 => 
                           n2805, QN => RAMDOUT1(5));
   U3294 : AOI221X1 port map( IN1 => RAM_12_5_port, IN2 => n2454, IN3 => 
                           RAM_13_5_port, IN4 => n3376, IN5 => n2848, QN => 
                           n2803);
   U3295 : AOI221X1 port map( IN1 => RAM_0_5_port, IN2 => n2172, IN3 => 
                           RAM_1_5_port, IN4 => n3390, IN5 => n2849, QN => 
                           n2804);
   U3296 : AOI221X2 port map( IN1 => RAM_4_5_port, IN2 => n3403, IN3 => 
                           RAM_5_5_port, IN4 => n3393, IN5 => n2850, QN => 
                           n2805);
   U3297 : NAND4X0 port map( IN1 => n2806, IN2 => n2808, IN3 => n2809, IN4 => 
                           n2807, QN => RAMDOUT1(125));
   U3298 : AOI221X1 port map( IN1 => RAM_8_125_port, IN2 => n3421, IN3 => 
                           RAM_9_125_port, IN4 => n3362, IN5 => n3331, QN => 
                           n2806);
   U3299 : AOI221X1 port map( IN1 => RAM_12_125_port, IN2 => n2459, IN3 => 
                           RAM_13_125_port, IN4 => n3375, IN5 => n3332, QN => 
                           n2807);
   U3300 : AOI221X1 port map( IN1 => RAM_0_125_port, IN2 => n2166, IN3 => 
                           RAM_1_125_port, IN4 => n3384, IN5 => n3333, QN => 
                           n2808);
   U3301 : AOI221X1 port map( IN1 => RAM_4_125_port, IN2 => n3406, IN3 => 
                           RAM_5_125_port, IN4 => n3398, IN5 => n3334, QN => 
                           n2809);
   U3302 : AO22X2 port map( IN1 => RAM_11_72_port, IN2 => n3462, IN3 => n2650, 
                           IN4 => RAM_10_72_port, Q => n3115);
   U3303 : AO22X2 port map( IN1 => RAM_11_62_port, IN2 => n3455, IN3 => 
                           RAM_10_62_port, IN4 => n2667, Q => n3075);
   U3304 : AO22X2 port map( IN1 => RAM_11_86_port, IN2 => n3458, IN3 => 
                           RAM_10_86_port, IN4 => n2666, Q => n3171);
   U3305 : AO22X2 port map( IN1 => RAM_11_9_port, IN2 => n2231, IN3 => n2665, 
                           IN4 => RAM_10_9_port, Q => n2863);
   U3306 : INVX0 port map( INP => n5616, ZN => n2810);
   U3307 : IBUFFX16 port map( INP => n2100, ZN => n5616);
   U3308 : AND2X4 port map( IN1 => n2821, IN2 => n2827, Q => n3344);
   U3309 : AND2X4 port map( IN1 => n2821, IN2 => n2827, Q => n3447);
   U3310 : AND2X4 port map( IN1 => n2825, IN2 => n2821, Q => n3347);
   U3311 : AND2X4 port map( IN1 => n2709, IN2 => n34, Q => n23);
   U3312 : AND2X4 port map( IN1 => n45, IN2 => n2709, Q => n37);
   U3313 : AND2X4 port map( IN1 => RAMADDR1(0), IN2 => RAMADDR1(1), Q => n2827)
                           ;
   U3314 : NAND4X0 port map( IN1 => n2811, IN2 => n2812, IN3 => n2813, IN4 => 
                           n2814, QN => RAMDOUT1(24));
   U3315 : AOI221X1 port map( IN1 => RAM_8_24_port, IN2 => n3420, IN3 => 
                           RAM_9_24_port, IN4 => n3365, IN5 => n2923, QN => 
                           n2811);
   U3316 : AOI221X1 port map( IN1 => RAM_12_24_port, IN2 => n2448, IN3 => 
                           RAM_13_24_port, IN4 => n3377, IN5 => n2924, QN => 
                           n2812);
   U3317 : AOI221X1 port map( IN1 => RAM_0_24_port, IN2 => n2162, IN3 => 
                           RAM_1_24_port, IN4 => n3386, IN5 => n2925, QN => 
                           n2813);
   U3318 : AOI221X1 port map( IN1 => RAM_4_24_port, IN2 => n3409, IN3 => 
                           RAM_5_24_port, IN4 => n3391, IN5 => n2926, QN => 
                           n2814);
   U3319 : NAND4X0 port map( IN1 => n2815, IN2 => n2816, IN3 => n2817, IN4 => 
                           n2818, QN => RAMDOUT1(113));
   U3320 : AOI221X1 port map( IN1 => RAM_8_113_port, IN2 => n3422, IN3 => 
                           RAM_9_113_port, IN4 => n3369, IN5 => n3283, QN => 
                           n2815);
   U3321 : AOI221X1 port map( IN1 => RAM_12_113_port, IN2 => n2455, IN3 => 
                           RAM_13_113_port, IN4 => n3375, IN5 => n3284, QN => 
                           n2816);
   U3322 : AOI221X1 port map( IN1 => RAM_0_113_port, IN2 => n2168, IN3 => 
                           RAM_1_113_port, IN4 => n3385, IN5 => n3285, QN => 
                           n2817);
   U3323 : AOI221X1 port map( IN1 => RAM_4_113_port, IN2 => n3402, IN3 => 
                           RAM_5_113_port, IN4 => n3398, IN5 => n3286, QN => 
                           n2818);
   U3324 : AO22X2 port map( IN1 => RAM_3_1_port, IN2 => n2548, IN3 => 
                           RAM_2_1_port, IN4 => n2629, Q => n2833);
   U3325 : AO22X2 port map( IN1 => RAM_3_73_port, IN2 => n2547, IN3 => n2099, 
                           IN4 => RAM_2_73_port, Q => n3121);
   U3326 : AO22X2 port map( IN1 => RAM_3_2_port, IN2 => n2469, IN3 => 
                           RAM_2_2_port, IN4 => n2644, Q => n2837);
   U3327 : AO22X2 port map( IN1 => RAM_3_52_port, IN2 => n2538, IN3 => 
                           RAM_2_52_port, IN4 => n2634, Q => n3037);
   U3328 : AO22X2 port map( IN1 => RAM_3_98_port, IN2 => n2399, IN3 => n2642, 
                           IN4 => RAM_2_98_port, Q => n3221);
   U3329 : AO22X2 port map( IN1 => RAM_3_11_port, IN2 => n2549, IN3 => 
                           RAM_2_11_port, IN4 => n2633, Q => n2873);
   U3330 : AO22X2 port map( IN1 => RAM_3_37_port, IN2 => n2545, IN3 => n2643, 
                           IN4 => RAM_2_37_port, Q => n2977);
   U3331 : AO22X2 port map( IN1 => RAM_3_21_port, IN2 => n2554, IN3 => 
                           RAM_2_21_port, IN4 => n2633, Q => n2913);
   U3332 : AO22X2 port map( IN1 => RAM_3_38_port, IN2 => n2552, IN3 => n2637, 
                           IN4 => RAM_2_38_port, Q => n2981);
   U3333 : AO22X2 port map( IN1 => RAM_3_62_port, IN2 => n2551, IN3 => 
                           RAM_2_62_port, IN4 => n2634, Q => n3077);
   U3334 : AO22X2 port map( IN1 => RAM_3_5_port, IN2 => n2551, IN3 => 
                           RAM_2_5_port, IN4 => n2627, Q => n2849);
   U3335 : AO22X2 port map( IN1 => RAM_3_58_port, IN2 => n2543, IN3 => 
                           RAM_2_58_port, IN4 => n2629, Q => n3061);
   U3336 : AO22X2 port map( IN1 => RAM_11_73_port, IN2 => n3450, IN3 => n2656, 
                           IN4 => RAM_10_73_port, Q => n3119);
   U3337 : AO22X2 port map( IN1 => RAM_11_102_port, IN2 => n3460, IN3 => 
                           RAM_10_102_port, IN4 => n2467, Q => n3235);
   U3338 : AO22X2 port map( IN1 => RAM_11_125_port, IN2 => n2466, IN3 => 
                           RAM_10_125_port, IN4 => n2467, Q => n3331);
   U3339 : AO22X2 port map( IN1 => RAM_11_38_port, IN2 => n2466, IN3 => 
                           RAM_10_38_port, IN4 => n2373, Q => n2979);
   U3340 : AO22X2 port map( IN1 => RAM_11_75_port, IN2 => n2498, IN3 => 
                           RAM_10_75_port, IN4 => n2655, Q => n3127);
   U3341 : AO22X2 port map( IN1 => RAM_11_33_port, IN2 => n3455, IN3 => 
                           RAM_10_33_port, IN4 => n2373, Q => n2959);
   U3342 : AO22X2 port map( IN1 => RAM_11_81_port, IN2 => n3458, IN3 => 
                           RAM_10_81_port, IN4 => n2664, Q => n3151);
   U3343 : AO22X2 port map( IN1 => RAM_11_68_port, IN2 => n3450, IN3 => 
                           RAM_10_68_port, IN4 => n2654, Q => n3099);
   U3344 : AO22X2 port map( IN1 => RAM_11_16_port, IN2 => n3460, IN3 => n2112, 
                           IN4 => RAM_10_16_port, Q => n2891);
   U3345 : AO22X2 port map( IN1 => RAM_11_60_port, IN2 => n3449, IN3 => n2664, 
                           IN4 => RAM_10_60_port, Q => n3067);
   U3346 : AO22X2 port map( IN1 => RAM_11_111_port, IN2 => n2231, IN3 => 
                           RAM_10_111_port, IN4 => n2653, Q => n3271);
   U3347 : AO22X2 port map( IN1 => RAM_11_123_port, IN2 => n2504, IN3 => n2652,
                           IN4 => RAM_10_123_port, Q => n3323);
   U3348 : AO22X2 port map( IN1 => RAM_11_127_port, IN2 => n3454, IN3 => 
                           RAM_10_127_port, IN4 => n2112, Q => n3341);
   U3349 : AO22X2 port map( IN1 => RAM_11_103_port, IN2 => n3449, IN3 => 
                           RAM_10_103_port, IN4 => n2657, Q => n3239);
   U3350 : AO22X2 port map( IN1 => RAM_11_121_port, IN2 => n3451, IN3 => 
                           RAM_10_121_port, IN4 => n2654, Q => n3315);
   U3351 : AO22X2 port map( IN1 => RAM_11_83_port, IN2 => n3449, IN3 => 
                           RAM_10_83_port, IN4 => n2655, Q => n3159);
   U3352 : AO22X2 port map( IN1 => RAM_11_78_port, IN2 => n3460, IN3 => 
                           RAM_10_78_port, IN4 => n2662, Q => n3139);
   U3353 : AO22X2 port map( IN1 => RAM_11_122_port, IN2 => n3450, IN3 => 
                           RAM_10_122_port, IN4 => n2461, Q => n3319);
   U3354 : AO22X2 port map( IN1 => RAM_7_54_port, IN2 => n2516, IN3 => 
                           RAM_6_54_port, IN4 => n2140, Q => n3046);
   U3355 : AO22X2 port map( IN1 => RAM_7_36_port, IN2 => n2515, IN3 => 
                           RAM_6_36_port, IN4 => n2137, Q => n2974);
   U3356 : AO22X2 port map( IN1 => RAM_7_102_port, IN2 => n2527, IN3 => 
                           RAM_6_102_port, IN4 => n2140, Q => n3238);
   U3357 : AO22X2 port map( IN1 => RAM_7_19_port, IN2 => n2521, IN3 => 
                           RAM_6_19_port, IN4 => n2136, Q => n2906);
   U3358 : AO22X2 port map( IN1 => RAM_7_60_port, IN2 => n2514, IN3 => 
                           RAM_6_60_port, IN4 => n2133, Q => n3070);
   U3359 : AO22X2 port map( IN1 => RAM_7_9_port, IN2 => n2394, IN3 => 
                           RAM_6_9_port, IN4 => n2152, Q => n2866);
   U3360 : AO22X2 port map( IN1 => RAM_7_83_port, IN2 => n2531, IN3 => 
                           RAM_6_83_port, IN4 => n2139, Q => n3162);
   U3361 : AO22X2 port map( IN1 => RAM_7_10_port, IN2 => n2523, IN3 => 
                           RAM_6_10_port, IN4 => n2137, Q => n2870);
   U3362 : AO22X2 port map( IN1 => RAM_7_116_port, IN2 => n2529, IN3 => 
                           RAM_6_116_port, IN4 => n2136, Q => n3298);
   U3363 : AO22X2 port map( IN1 => n2501, IN2 => RAM_11_85_port, IN3 => 
                           RAM_10_85_port, IN4 => n2467, Q => n3167);
   U3364 : AO22X2 port map( IN1 => RAM_11_109_port, IN2 => n2466, IN3 => 
                           RAM_10_109_port, IN4 => n2661, Q => n3263);
   U3365 : AO22X2 port map( IN1 => RAM_11_5_port, IN2 => n3455, IN3 => 
                           RAM_10_5_port, IN4 => n2667, Q => n2847);
   U3366 : AO22X2 port map( IN1 => RAM_11_27_port, IN2 => n2231, IN3 => n2651, 
                           IN4 => RAM_10_27_port, Q => n2935);
   U3367 : AO22X2 port map( IN1 => RAM_11_14_port, IN2 => n3458, IN3 => 
                           RAM_10_14_port, IN4 => n2658, Q => n2883);
   U3368 : AO22X2 port map( IN1 => RAM_11_98_port, IN2 => n3460, IN3 => n2373, 
                           IN4 => RAM_10_98_port, Q => n3219);
   U3369 : AO22X2 port map( IN1 => RAM_11_115_port, IN2 => n3454, IN3 => 
                           RAM_10_115_port, IN4 => n2652, Q => n3291);
   U3370 : AO22X2 port map( IN1 => RAM_11_104_port, IN2 => n2231, IN3 => n2665,
                           IN4 => RAM_10_104_port, Q => n3243);
   U3371 : AO22X2 port map( IN1 => RAM_11_112_port, IN2 => n3458, IN3 => n2665,
                           IN4 => RAM_10_112_port, Q => n3275);
   U3372 : AO22X2 port map( IN1 => RAM_11_71_port, IN2 => n3454, IN3 => n2652, 
                           IN4 => RAM_10_71_port, Q => n3111);
   U3373 : AO22X2 port map( IN1 => RAM_11_94_port, IN2 => n3461, IN3 => n2480, 
                           IN4 => RAM_10_94_port, Q => n3203);
   U3374 : AO22X2 port map( IN1 => RAM_15_108_port, IN2 => n3440, IN3 => 
                           RAM_14_108_port, IN4 => n2326, Q => n3260);
   U3375 : AO22X2 port map( IN1 => RAM_15_40_port, IN2 => n3446, IN3 => 
                           RAM_14_40_port, IN4 => n2328, Q => n2988);
   U3376 : AO22X2 port map( IN1 => RAM_15_77_port, IN2 => n3441, IN3 => 
                           RAM_14_77_port, IN4 => n2333, Q => n3136);
   U3377 : AO22X2 port map( IN1 => RAM_15_11_port, IN2 => n3440, IN3 => 
                           RAM_14_11_port, IN4 => n2329, Q => n2872);
   U3378 : AO22X2 port map( IN1 => RAM_15_41_port, IN2 => n3439, IN3 => 
                           RAM_14_41_port, IN4 => n2326, Q => n2992);
   U3379 : AO22X2 port map( IN1 => RAM_15_98_port, IN2 => n3441, IN3 => 
                           RAM_14_98_port, IN4 => n2320, Q => n3220);
   U3380 : AO22X2 port map( IN1 => RAM_15_127_port, IN2 => n3433, IN3 => 
                           RAM_14_127_port, IN4 => n2339, Q => n3345);
   U3381 : AO22X2 port map( IN1 => RAM_15_103_port, IN2 => n3445, IN3 => 
                           RAM_14_103_port, IN4 => n2329, Q => n3240);
   U3382 : AO22X2 port map( IN1 => RAM_15_28_port, IN2 => n3437, IN3 => 
                           RAM_14_28_port, IN4 => n2331, Q => n2940);
   U3383 : AO22X2 port map( IN1 => RAM_15_102_port, IN2 => n3436, IN3 => 
                           RAM_14_102_port, IN4 => n2327, Q => n3236);
   U3384 : AO22X2 port map( IN1 => RAM_15_119_port, IN2 => n3434, IN3 => 
                           RAM_14_119_port, IN4 => n2325, Q => n3308);
   U3385 : AO22X2 port map( IN1 => RAM_15_24_port, IN2 => n3437, IN3 => 
                           RAM_14_24_port, IN4 => n2328, Q => n2924);
   U3386 : AO22X2 port map( IN1 => RAM_15_58_port, IN2 => n3445, IN3 => 
                           RAM_14_58_port, IN4 => n2333, Q => n3060);
   U3387 : AO22X2 port map( IN1 => RAM_15_101_port, IN2 => n3439, IN3 => 
                           RAM_14_101_port, IN4 => n2335, Q => n3232);
   U3388 : AO22X2 port map( IN1 => RAM_15_99_port, IN2 => n3446, IN3 => 
                           RAM_14_99_port, IN4 => n2330, Q => n3224);
   U3389 : NBUFFX2 port map( INP => n4499, Z => n4605);
   U3390 : NBUFFX2 port map( INP => n4504, Z => n4649);
   U3391 : NBUFFX2 port map( INP => n4489, Z => n4517);
   U3392 : NBUFFX2 port map( INP => n4499, Z => n4614);
   U3393 : NBUFFX2 port map( INP => n4504, Z => n4658);
   U3394 : NBUFFX2 port map( INP => n4489, Z => n4526);
   U3395 : NBUFFX2 port map( INP => n4494, Z => n4570);
   U3396 : NBUFFX2 port map( INP => n4494, Z => n4561);
   U3397 : NBUFFX2 port map( INP => n4489, Z => n4525);
   U3398 : NBUFFX2 port map( INP => n4489, Z => n4524);
   U3399 : NBUFFX2 port map( INP => n4504, Z => n4657);
   U3400 : NBUFFX2 port map( INP => n4504, Z => n4656);
   U3401 : NBUFFX2 port map( INP => n4499, Z => n4613);
   U3402 : NBUFFX2 port map( INP => n4499, Z => n4612);
   U3403 : NBUFFX2 port map( INP => n4495, Z => n4581);
   U3404 : NBUFFX2 port map( INP => n4495, Z => n4572);
   U3405 : NBUFFX2 port map( INP => n4505, Z => n4660);
   U3406 : NBUFFX2 port map( INP => n4505, Z => n4669);
   U3407 : NBUFFX2 port map( INP => n4505, Z => n4668);
   U3408 : NBUFFX2 port map( INP => n4505, Z => n4667);
   U3409 : NBUFFX2 port map( INP => n4507, Z => n4679);
   U3410 : NBUFFX2 port map( INP => n4502, Z => n4635);
   U3411 : NBUFFX2 port map( INP => n4507, Z => n4678);
   U3412 : NBUFFX2 port map( INP => n4502, Z => n4634);
   U3413 : NBUFFX2 port map( INP => n4492, Z => n4547);
   U3414 : NBUFFX2 port map( INP => n4492, Z => n4546);
   U3415 : NBUFFX2 port map( INP => n4497, Z => n4583);
   U3416 : NBUFFX2 port map( INP => n4497, Z => n4592);
   U3417 : NBUFFX2 port map( INP => n4498, Z => n4594);
   U3418 : NBUFFX2 port map( INP => n4498, Z => n4603);
   U3419 : NBUFFX2 port map( INP => n4508, Z => n4691);
   U3420 : NBUFFX2 port map( INP => n4508, Z => n4682);
   U3421 : NBUFFX2 port map( INP => n4508, Z => n4690);
   U3422 : NBUFFX2 port map( INP => n4508, Z => n4689);
   U3423 : NBUFFX2 port map( INP => n4493, Z => n4558);
   U3424 : NBUFFX2 port map( INP => n4493, Z => n4557);
   U3425 : NBUFFX2 port map( INP => n4503, Z => n4646);
   U3426 : NBUFFX2 port map( INP => n4503, Z => n4645);
   U3427 : NBUFFX2 port map( INP => n4490, Z => n4528);
   U3428 : NBUFFX2 port map( INP => n4500, Z => n4616);
   U3429 : NBUFFX2 port map( INP => n4490, Z => n4537);
   U3430 : NBUFFX2 port map( INP => n4500, Z => n4625);
   U3431 : NBUFFX2 port map( INP => n4500, Z => n4624);
   U3432 : NBUFFX2 port map( INP => n4500, Z => n4623);
   U3433 : NBUFFX2 port map( INP => n4490, Z => n4536);
   U3434 : NBUFFX2 port map( INP => n4490, Z => n4535);
   U3435 : INVX0 port map( INP => n5047, ZN => n5045);
   U3436 : INVX0 port map( INP => n5047, ZN => n5044);
   U3437 : INVX0 port map( INP => n5047, ZN => n5043);
   U3438 : INVX0 port map( INP => n5047, ZN => n5042);
   U3439 : INVX0 port map( INP => n5048, ZN => n5041);
   U3440 : INVX0 port map( INP => n5048, ZN => n5040);
   U3441 : INVX0 port map( INP => n5048, ZN => n5039);
   U3442 : INVX0 port map( INP => n5048, ZN => n5038);
   U3443 : INVX0 port map( INP => n5048, ZN => n5037);
   U3444 : INVX0 port map( INP => n5048, ZN => n5036);
   U3445 : INVX0 port map( INP => n5214, ZN => n5212);
   U3446 : INVX0 port map( INP => n5214, ZN => n5211);
   U3447 : INVX0 port map( INP => n5214, ZN => n5210);
   U3448 : INVX0 port map( INP => n5214, ZN => n5209);
   U3449 : INVX0 port map( INP => n5215, ZN => n5208);
   U3450 : INVX0 port map( INP => n5215, ZN => n5207);
   U3451 : INVX0 port map( INP => n5215, ZN => n5206);
   U3452 : INVX0 port map( INP => n5215, ZN => n5205);
   U3453 : INVX0 port map( INP => n5215, ZN => n5204);
   U3454 : INVX0 port map( INP => n5215, ZN => n5203);
   U3455 : INVX0 port map( INP => n5549, ZN => n5541);
   U3456 : INVX0 port map( INP => n5549, ZN => n5540);
   U3457 : INVX0 port map( INP => n5549, ZN => n5539);
   U3458 : INVX0 port map( INP => n5549, ZN => n5538);
   U3459 : INVX0 port map( INP => n5549, ZN => n5537);
   U3460 : INVX0 port map( INP => n5382, ZN => n5380);
   U3461 : INVX0 port map( INP => n5382, ZN => n5379);
   U3462 : INVX0 port map( INP => n5382, ZN => n5378);
   U3463 : INVX0 port map( INP => n5382, ZN => n5377);
   U3464 : INVX0 port map( INP => n5383, ZN => n5376);
   U3465 : INVX0 port map( INP => n5383, ZN => n5375);
   U3466 : INVX0 port map( INP => n5383, ZN => n5374);
   U3467 : INVX0 port map( INP => n5383, ZN => n5373);
   U3468 : INVX0 port map( INP => n5383, ZN => n5372);
   U3469 : INVX0 port map( INP => n5383, ZN => n5371);
   U3470 : INVX0 port map( INP => n5548, ZN => n5545);
   U3471 : INVX0 port map( INP => n5548, ZN => n5544);
   U3472 : INVX0 port map( INP => n5548, ZN => n5543);
   U3473 : INVX0 port map( INP => n5549, ZN => n5542);
   U3474 : INVX0 port map( INP => n5047, ZN => n5046);
   U3475 : INVX0 port map( INP => n5214, ZN => n5213);
   U3476 : INVX0 port map( INP => n5382, ZN => n5381);
   U3477 : INVX0 port map( INP => n5548, ZN => n5547);
   U3478 : INVX0 port map( INP => n5030, ZN => n5049);
   U3479 : INVX0 port map( INP => n5030, ZN => n5050);
   U3480 : INVX0 port map( INP => n5030, ZN => n5051);
   U3481 : INVX0 port map( INP => n5030, ZN => n5052);
   U3482 : INVX0 port map( INP => n5030, ZN => n5053);
   U3483 : INVX0 port map( INP => n5031, ZN => n5054);
   U3484 : INVX0 port map( INP => n5031, ZN => n5055);
   U3485 : INVX0 port map( INP => n5031, ZN => n5056);
   U3486 : INVX0 port map( INP => n5031, ZN => n5057);
   U3487 : INVX0 port map( INP => n5031, ZN => n5058);
   U3488 : INVX0 port map( INP => n5032, ZN => n5059);
   U3489 : INVX0 port map( INP => n5032, ZN => n5060);
   U3490 : INVX0 port map( INP => n5032, ZN => n5061);
   U3491 : INVX0 port map( INP => n5032, ZN => n5062);
   U3492 : INVX0 port map( INP => n5032, ZN => n5063);
   U3493 : INVX0 port map( INP => n5033, ZN => n5064);
   U3494 : INVX0 port map( INP => n5033, ZN => n5065);
   U3495 : INVX0 port map( INP => n5033, ZN => n5066);
   U3496 : INVX0 port map( INP => n5033, ZN => n5067);
   U3497 : INVX0 port map( INP => n5033, ZN => n5068);
   U3498 : INVX0 port map( INP => n5197, ZN => n5216);
   U3499 : INVX0 port map( INP => n5197, ZN => n5217);
   U3500 : INVX0 port map( INP => n5197, ZN => n5218);
   U3501 : INVX0 port map( INP => n5197, ZN => n5219);
   U3502 : INVX0 port map( INP => n5197, ZN => n5220);
   U3503 : INVX0 port map( INP => n5198, ZN => n5221);
   U3504 : INVX0 port map( INP => n5198, ZN => n5222);
   U3505 : INVX0 port map( INP => n5198, ZN => n5223);
   U3506 : INVX0 port map( INP => n5198, ZN => n5224);
   U3507 : INVX0 port map( INP => n5198, ZN => n5225);
   U3508 : INVX0 port map( INP => n5199, ZN => n5226);
   U3509 : INVX0 port map( INP => n5199, ZN => n5227);
   U3510 : INVX0 port map( INP => n5199, ZN => n5228);
   U3511 : INVX0 port map( INP => n5199, ZN => n5229);
   U3512 : INVX0 port map( INP => n5199, ZN => n5230);
   U3513 : INVX0 port map( INP => n5200, ZN => n5231);
   U3514 : INVX0 port map( INP => n5200, ZN => n5232);
   U3515 : INVX0 port map( INP => n5200, ZN => n5233);
   U3516 : INVX0 port map( INP => n5200, ZN => n5234);
   U3517 : INVX0 port map( INP => n5200, ZN => n5235);
   U3518 : INVX0 port map( INP => n5548, ZN => n5546);
   U3519 : INVX0 port map( INP => n5532, ZN => n5559);
   U3520 : INVX0 port map( INP => n5533, ZN => n5560);
   U3521 : INVX0 port map( INP => n5532, ZN => n5558);
   U3522 : INVX0 port map( INP => n5034, ZN => n5069);
   U3523 : INVX0 port map( INP => n5034, ZN => n5070);
   U3524 : INVX0 port map( INP => n5201, ZN => n5236);
   U3525 : INVX0 port map( INP => n5201, ZN => n5237);
   U3526 : INVX0 port map( INP => n5531, ZN => n5550);
   U3527 : INVX0 port map( INP => n5531, ZN => n5551);
   U3528 : INVX0 port map( INP => n5531, ZN => n5552);
   U3529 : INVX0 port map( INP => n5531, ZN => n5553);
   U3530 : INVX0 port map( INP => n5531, ZN => n5554);
   U3531 : INVX0 port map( INP => n5532, ZN => n5555);
   U3532 : INVX0 port map( INP => n5532, ZN => n5556);
   U3533 : INVX0 port map( INP => n5532, ZN => n5557);
   U3534 : INVX0 port map( INP => n5533, ZN => n5561);
   U3535 : INVX0 port map( INP => n5533, ZN => n5562);
   U3536 : INVX0 port map( INP => n5533, ZN => n5563);
   U3537 : INVX0 port map( INP => n5533, ZN => n5564);
   U3538 : INVX0 port map( INP => n5534, ZN => n5565);
   U3539 : INVX0 port map( INP => n5534, ZN => n5566);
   U3540 : INVX0 port map( INP => n5534, ZN => n5567);
   U3541 : INVX0 port map( INP => n5534, ZN => n5568);
   U3542 : INVX0 port map( INP => n5534, ZN => n5569);
   U3543 : INVX0 port map( INP => n5365, ZN => n5384);
   U3544 : INVX0 port map( INP => n5365, ZN => n5385);
   U3545 : INVX0 port map( INP => n5365, ZN => n5386);
   U3546 : INVX0 port map( INP => n5365, ZN => n5387);
   U3547 : INVX0 port map( INP => n5366, ZN => n5388);
   U3548 : INVX0 port map( INP => n5366, ZN => n5389);
   U3549 : INVX0 port map( INP => n5366, ZN => n5390);
   U3550 : INVX0 port map( INP => n5366, ZN => n5391);
   U3551 : INVX0 port map( INP => n5366, ZN => n5392);
   U3552 : INVX0 port map( INP => n5367, ZN => n5393);
   U3553 : INVX0 port map( INP => n5367, ZN => n5394);
   U3554 : INVX0 port map( INP => n5367, ZN => n5395);
   U3555 : INVX0 port map( INP => n5367, ZN => n5396);
   U3556 : INVX0 port map( INP => n5367, ZN => n5397);
   U3557 : INVX0 port map( INP => n5368, ZN => n5398);
   U3558 : INVX0 port map( INP => n5368, ZN => n5399);
   U3559 : INVX0 port map( INP => n5368, ZN => n5400);
   U3560 : INVX0 port map( INP => n5368, ZN => n5401);
   U3561 : INVX0 port map( INP => n5368, ZN => n5402);
   U3562 : INVX0 port map( INP => n5535, ZN => n5570);
   U3563 : INVX0 port map( INP => n5535, ZN => n5571);
   U3564 : INVX0 port map( INP => n5369, ZN => n5403);
   U3565 : INVX0 port map( INP => n5369, ZN => n5404);
   U3566 : INVX0 port map( INP => n5034, ZN => n5071);
   U3567 : INVX0 port map( INP => n5201, ZN => n5238);
   U3568 : INVX0 port map( INP => n5535, ZN => n5572);
   U3569 : INVX0 port map( INP => n5369, ZN => n5405);
   U3570 : INVX0 port map( INP => n5591, ZN => n5583);
   U3571 : INVX0 port map( INP => n5590, ZN => n5588);
   U3572 : INVX0 port map( INP => n5590, ZN => n5587);
   U3573 : INVX0 port map( INP => n5590, ZN => n5586);
   U3574 : INVX0 port map( INP => n5590, ZN => n5585);
   U3575 : INVX0 port map( INP => n5591, ZN => n5582);
   U3576 : INVX0 port map( INP => n5591, ZN => n5581);
   U3577 : INVX0 port map( INP => n5591, ZN => n5580);
   U3578 : INVX0 port map( INP => n5590, ZN => n5579);
   U3579 : INVX0 port map( INP => n5506, ZN => n5504);
   U3580 : INVX0 port map( INP => n5506, ZN => n5503);
   U3581 : INVX0 port map( INP => n5506, ZN => n5502);
   U3582 : INVX0 port map( INP => n5506, ZN => n5501);
   U3583 : INVX0 port map( INP => n5507, ZN => n5500);
   U3584 : INVX0 port map( INP => n5507, ZN => n5499);
   U3585 : INVX0 port map( INP => n5507, ZN => n5498);
   U3586 : INVX0 port map( INP => n5507, ZN => n5497);
   U3587 : INVX0 port map( INP => n5507, ZN => n5496);
   U3588 : INVX0 port map( INP => n5507, ZN => n5495);
   U3589 : INVX0 port map( INP => n5464, ZN => n5462);
   U3590 : INVX0 port map( INP => n5464, ZN => n5461);
   U3591 : INVX0 port map( INP => n5464, ZN => n5460);
   U3592 : INVX0 port map( INP => n5464, ZN => n5459);
   U3593 : INVX0 port map( INP => n5465, ZN => n5458);
   U3594 : INVX0 port map( INP => n5465, ZN => n5457);
   U3595 : INVX0 port map( INP => n5465, ZN => n5456);
   U3596 : INVX0 port map( INP => n5465, ZN => n5455);
   U3597 : INVX0 port map( INP => n5465, ZN => n5454);
   U3598 : INVX0 port map( INP => n5465, ZN => n5453);
   U3599 : INVX0 port map( INP => n5172, ZN => n5170);
   U3600 : INVX0 port map( INP => n5172, ZN => n5169);
   U3601 : INVX0 port map( INP => n5172, ZN => n5168);
   U3602 : INVX0 port map( INP => n5172, ZN => n5167);
   U3603 : INVX0 port map( INP => n5173, ZN => n5166);
   U3604 : INVX0 port map( INP => n5173, ZN => n5165);
   U3605 : INVX0 port map( INP => n5173, ZN => n5164);
   U3606 : INVX0 port map( INP => n5173, ZN => n5163);
   U3607 : INVX0 port map( INP => n5173, ZN => n5162);
   U3608 : INVX0 port map( INP => n5130, ZN => n5128);
   U3609 : INVX0 port map( INP => n5130, ZN => n5127);
   U3610 : INVX0 port map( INP => n5130, ZN => n5126);
   U3611 : INVX0 port map( INP => n5130, ZN => n5125);
   U3612 : INVX0 port map( INP => n5131, ZN => n5124);
   U3613 : INVX0 port map( INP => n5131, ZN => n5123);
   U3614 : INVX0 port map( INP => n5131, ZN => n5122);
   U3615 : INVX0 port map( INP => n5131, ZN => n5121);
   U3616 : INVX0 port map( INP => n5131, ZN => n5120);
   U3617 : INVX0 port map( INP => n5173, ZN => n5161);
   U3618 : INVX0 port map( INP => n5131, ZN => n5119);
   U3619 : INVX0 port map( INP => n5340, ZN => n5338);
   U3620 : INVX0 port map( INP => n5340, ZN => n5337);
   U3621 : INVX0 port map( INP => n5340, ZN => n5336);
   U3622 : INVX0 port map( INP => n5340, ZN => n5335);
   U3623 : INVX0 port map( INP => n5340, ZN => n5329);
   U3624 : INVX0 port map( INP => n5423, ZN => n5421);
   U3625 : INVX0 port map( INP => n5423, ZN => n5420);
   U3626 : INVX0 port map( INP => n5423, ZN => n5419);
   U3627 : INVX0 port map( INP => n5423, ZN => n5418);
   U3628 : INVX0 port map( INP => n5423, ZN => n5412);
   U3629 : INVX0 port map( INP => n5005, ZN => n5003);
   U3630 : INVX0 port map( INP => n5005, ZN => n5002);
   U3631 : INVX0 port map( INP => n5005, ZN => n5001);
   U3632 : INVX0 port map( INP => n5005, ZN => n5000);
   U3633 : INVX0 port map( INP => n5006, ZN => n4999);
   U3634 : INVX0 port map( INP => n5006, ZN => n4998);
   U3635 : INVX0 port map( INP => n5006, ZN => n4997);
   U3636 : INVX0 port map( INP => n5006, ZN => n4996);
   U3637 : INVX0 port map( INP => n5006, ZN => n4995);
   U3638 : INVX0 port map( INP => n5005, ZN => n4994);
   U3639 : INVX0 port map( INP => n5089, ZN => n5087);
   U3640 : INVX0 port map( INP => n5089, ZN => n5086);
   U3641 : INVX0 port map( INP => n5089, ZN => n5085);
   U3642 : INVX0 port map( INP => n5089, ZN => n5084);
   U3643 : INVX0 port map( INP => n5090, ZN => n5083);
   U3644 : INVX0 port map( INP => n5090, ZN => n5082);
   U3645 : INVX0 port map( INP => n5090, ZN => n5081);
   U3646 : INVX0 port map( INP => n5090, ZN => n5080);
   U3647 : INVX0 port map( INP => n5090, ZN => n5079);
   U3648 : INVX0 port map( INP => n5090, ZN => n5078);
   U3649 : INVX0 port map( INP => n5256, ZN => n5254);
   U3650 : INVX0 port map( INP => n5256, ZN => n5253);
   U3651 : INVX0 port map( INP => n5256, ZN => n5252);
   U3652 : INVX0 port map( INP => n5256, ZN => n5251);
   U3653 : INVX0 port map( INP => n5257, ZN => n5250);
   U3654 : INVX0 port map( INP => n5257, ZN => n5249);
   U3655 : INVX0 port map( INP => n5257, ZN => n5248);
   U3656 : INVX0 port map( INP => n5257, ZN => n5247);
   U3657 : INVX0 port map( INP => n5257, ZN => n5246);
   U3658 : INVX0 port map( INP => n5257, ZN => n5245);
   U3659 : INVX0 port map( INP => n4963, ZN => n4961);
   U3660 : INVX0 port map( INP => n4963, ZN => n4960);
   U3661 : INVX0 port map( INP => n4963, ZN => n4959);
   U3662 : INVX0 port map( INP => n4963, ZN => n4958);
   U3663 : INVX0 port map( INP => n4964, ZN => n4957);
   U3664 : INVX0 port map( INP => n4964, ZN => n4956);
   U3665 : INVX0 port map( INP => n4964, ZN => n4955);
   U3666 : INVX0 port map( INP => n4964, ZN => n4954);
   U3667 : INVX0 port map( INP => n4964, ZN => n4953);
   U3668 : INVX0 port map( INP => n4963, ZN => n4952);
   U3669 : INVX0 port map( INP => n5424, ZN => n5416);
   U3670 : INVX0 port map( INP => n5424, ZN => n5415);
   U3671 : INVX0 port map( INP => n5424, ZN => n5414);
   U3672 : INVX0 port map( INP => n5424, ZN => n5413);
   U3673 : INVX0 port map( INP => n5341, ZN => n5333);
   U3674 : INVX0 port map( INP => n5341, ZN => n5332);
   U3675 : INVX0 port map( INP => n5341, ZN => n5331);
   U3676 : INVX0 port map( INP => n5341, ZN => n5330);
   U3677 : INVX0 port map( INP => n5590, ZN => n5589);
   U3678 : INVX0 port map( INP => n5506, ZN => n5505);
   U3679 : INVX0 port map( INP => n5464, ZN => n5463);
   U3680 : INVX0 port map( INP => n5172, ZN => n5171);
   U3681 : INVX0 port map( INP => n5130, ZN => n5129);
   U3682 : INVX0 port map( INP => n5340, ZN => n5339);
   U3683 : INVX0 port map( INP => n5423, ZN => n5422);
   U3684 : INVX0 port map( INP => n5005, ZN => n5004);
   U3685 : INVX0 port map( INP => n5089, ZN => n5088);
   U3686 : INVX0 port map( INP => n5256, ZN => n5255);
   U3687 : INVX0 port map( INP => n43, ZN => n5048);
   U3688 : INVX0 port map( INP => n38, ZN => n5215);
   U3689 : INVX0 port map( INP => n43, ZN => n5047);
   U3690 : INVX0 port map( INP => n38, ZN => n5214);
   U3691 : INVX0 port map( INP => n5424, ZN => n5417);
   U3692 : INVX0 port map( INP => n5591, ZN => n5584);
   U3693 : INVX0 port map( INP => n5298, ZN => n5296);
   U3694 : INVX0 port map( INP => n5298, ZN => n5295);
   U3695 : INVX0 port map( INP => n5298, ZN => n5294);
   U3696 : INVX0 port map( INP => n5298, ZN => n5293);
   U3697 : INVX0 port map( INP => n5299, ZN => n5292);
   U3698 : INVX0 port map( INP => n5299, ZN => n5291);
   U3699 : INVX0 port map( INP => n5299, ZN => n5290);
   U3700 : INVX0 port map( INP => n5299, ZN => n5289);
   U3701 : INVX0 port map( INP => n5299, ZN => n5288);
   U3702 : INVX0 port map( INP => n5299, ZN => n5287);
   U3703 : INVX0 port map( INP => n4963, ZN => n4962);
   U3704 : INVX0 port map( INP => n5298, ZN => n5297);
   U3705 : INVX0 port map( INP => n24, ZN => n5549);
   U3706 : INVX0 port map( INP => n31, ZN => n5383);
   U3707 : INVX0 port map( INP => n31, ZN => n5382);
   U3708 : INVX0 port map( INP => n5035, ZN => n5030);
   U3709 : INVX0 port map( INP => n5035, ZN => n5031);
   U3710 : INVX0 port map( INP => n5035, ZN => n5032);
   U3711 : INVX0 port map( INP => n5035, ZN => n5033);
   U3712 : INVX0 port map( INP => n5202, ZN => n5197);
   U3713 : INVX0 port map( INP => n5202, ZN => n5198);
   U3714 : INVX0 port map( INP => n5202, ZN => n5199);
   U3715 : INVX0 port map( INP => n5202, ZN => n5200);
   U3716 : INVX0 port map( INP => n5574, ZN => n5600);
   U3717 : INVX0 port map( INP => n5323, ZN => n5342);
   U3718 : INVX0 port map( INP => n5323, ZN => n5343);
   U3719 : INVX0 port map( INP => n5323, ZN => n5344);
   U3720 : INVX0 port map( INP => n5323, ZN => n5345);
   U3721 : INVX0 port map( INP => n5323, ZN => n5346);
   U3722 : INVX0 port map( INP => n5324, ZN => n5347);
   U3723 : INVX0 port map( INP => n5324, ZN => n5348);
   U3724 : INVX0 port map( INP => n5324, ZN => n5349);
   U3725 : INVX0 port map( INP => n5324, ZN => n5350);
   U3726 : INVX0 port map( INP => n5324, ZN => n5351);
   U3727 : INVX0 port map( INP => n5325, ZN => n5352);
   U3728 : INVX0 port map( INP => n5325, ZN => n5353);
   U3729 : INVX0 port map( INP => n5325, ZN => n5354);
   U3730 : INVX0 port map( INP => n5325, ZN => n5355);
   U3731 : INVX0 port map( INP => n5325, ZN => n5356);
   U3732 : INVX0 port map( INP => n5326, ZN => n5357);
   U3733 : INVX0 port map( INP => n5326, ZN => n5358);
   U3734 : INVX0 port map( INP => n5326, ZN => n5359);
   U3735 : INVX0 port map( INP => n5326, ZN => n5360);
   U3736 : INVX0 port map( INP => n5326, ZN => n5361);
   U3737 : INVX0 port map( INP => n5406, ZN => n5425);
   U3738 : INVX0 port map( INP => n5406, ZN => n5426);
   U3739 : INVX0 port map( INP => n5406, ZN => n5427);
   U3740 : INVX0 port map( INP => n5406, ZN => n5428);
   U3741 : INVX0 port map( INP => n5407, ZN => n5429);
   U3742 : INVX0 port map( INP => n5407, ZN => n5430);
   U3743 : INVX0 port map( INP => n5407, ZN => n5431);
   U3744 : INVX0 port map( INP => n5407, ZN => n5432);
   U3745 : INVX0 port map( INP => n5407, ZN => n5433);
   U3746 : INVX0 port map( INP => n5408, ZN => n5434);
   U3747 : INVX0 port map( INP => n5408, ZN => n5435);
   U3748 : INVX0 port map( INP => n5408, ZN => n5436);
   U3749 : INVX0 port map( INP => n5408, ZN => n5437);
   U3750 : INVX0 port map( INP => n5408, ZN => n5438);
   U3751 : INVX0 port map( INP => n5409, ZN => n5439);
   U3752 : INVX0 port map( INP => n5409, ZN => n5440);
   U3753 : INVX0 port map( INP => n5409, ZN => n5441);
   U3754 : INVX0 port map( INP => n5409, ZN => n5442);
   U3755 : INVX0 port map( INP => n5409, ZN => n5443);
   U3756 : INVX0 port map( INP => n5327, ZN => n5362);
   U3757 : INVX0 port map( INP => n5327, ZN => n5363);
   U3758 : INVX0 port map( INP => n5410, ZN => n5444);
   U3759 : INVX0 port map( INP => n5410, ZN => n5445);
   U3760 : INVX0 port map( INP => n5489, ZN => n5508);
   U3761 : INVX0 port map( INP => n5489, ZN => n5509);
   U3762 : INVX0 port map( INP => n5489, ZN => n5510);
   U3763 : INVX0 port map( INP => n5489, ZN => n5511);
   U3764 : INVX0 port map( INP => n5489, ZN => n5512);
   U3765 : INVX0 port map( INP => n5490, ZN => n5513);
   U3766 : INVX0 port map( INP => n5490, ZN => n5514);
   U3767 : INVX0 port map( INP => n5490, ZN => n5515);
   U3768 : INVX0 port map( INP => n5490, ZN => n5516);
   U3769 : INVX0 port map( INP => n5490, ZN => n5517);
   U3770 : INVX0 port map( INP => n5491, ZN => n5518);
   U3771 : INVX0 port map( INP => n5491, ZN => n5519);
   U3772 : INVX0 port map( INP => n5491, ZN => n5520);
   U3773 : INVX0 port map( INP => n5491, ZN => n5521);
   U3774 : INVX0 port map( INP => n5491, ZN => n5522);
   U3775 : INVX0 port map( INP => n5492, ZN => n5523);
   U3776 : INVX0 port map( INP => n5492, ZN => n5524);
   U3777 : INVX0 port map( INP => n5492, ZN => n5525);
   U3778 : INVX0 port map( INP => n5492, ZN => n5526);
   U3779 : INVX0 port map( INP => n5492, ZN => n5527);
   U3780 : INVX0 port map( INP => n5447, ZN => n5466);
   U3781 : INVX0 port map( INP => n5447, ZN => n5467);
   U3782 : INVX0 port map( INP => n5447, ZN => n5468);
   U3783 : INVX0 port map( INP => n5447, ZN => n5469);
   U3784 : INVX0 port map( INP => n5447, ZN => n5470);
   U3785 : INVX0 port map( INP => n5448, ZN => n5471);
   U3786 : INVX0 port map( INP => n5448, ZN => n5472);
   U3787 : INVX0 port map( INP => n5448, ZN => n5473);
   U3788 : INVX0 port map( INP => n5448, ZN => n5474);
   U3789 : INVX0 port map( INP => n5448, ZN => n5475);
   U3790 : INVX0 port map( INP => n5449, ZN => n5476);
   U3791 : INVX0 port map( INP => n5449, ZN => n5477);
   U3792 : INVX0 port map( INP => n5449, ZN => n5478);
   U3793 : INVX0 port map( INP => n5449, ZN => n5479);
   U3794 : INVX0 port map( INP => n5449, ZN => n5480);
   U3795 : INVX0 port map( INP => n5450, ZN => n5481);
   U3796 : INVX0 port map( INP => n5450, ZN => n5482);
   U3797 : INVX0 port map( INP => n5450, ZN => n5483);
   U3798 : INVX0 port map( INP => n5450, ZN => n5484);
   U3799 : INVX0 port map( INP => n5450, ZN => n5485);
   U3800 : INVX0 port map( INP => n5155, ZN => n5174);
   U3801 : INVX0 port map( INP => n5155, ZN => n5175);
   U3802 : INVX0 port map( INP => n5155, ZN => n5176);
   U3803 : INVX0 port map( INP => n5155, ZN => n5177);
   U3804 : INVX0 port map( INP => n5155, ZN => n5178);
   U3805 : INVX0 port map( INP => n5156, ZN => n5179);
   U3806 : INVX0 port map( INP => n5156, ZN => n5180);
   U3807 : INVX0 port map( INP => n5156, ZN => n5181);
   U3808 : INVX0 port map( INP => n5156, ZN => n5182);
   U3809 : INVX0 port map( INP => n5156, ZN => n5183);
   U3810 : INVX0 port map( INP => n5157, ZN => n5184);
   U3811 : INVX0 port map( INP => n5157, ZN => n5185);
   U3812 : INVX0 port map( INP => n5157, ZN => n5186);
   U3813 : INVX0 port map( INP => n5157, ZN => n5187);
   U3814 : INVX0 port map( INP => n5157, ZN => n5188);
   U3815 : INVX0 port map( INP => n5158, ZN => n5189);
   U3816 : INVX0 port map( INP => n5158, ZN => n5190);
   U3817 : INVX0 port map( INP => n5158, ZN => n5191);
   U3818 : INVX0 port map( INP => n5158, ZN => n5192);
   U3819 : INVX0 port map( INP => n5158, ZN => n5193);
   U3820 : INVX0 port map( INP => n5113, ZN => n5132);
   U3821 : INVX0 port map( INP => n5113, ZN => n5133);
   U3822 : INVX0 port map( INP => n5113, ZN => n5134);
   U3823 : INVX0 port map( INP => n5113, ZN => n5135);
   U3824 : INVX0 port map( INP => n5113, ZN => n5136);
   U3825 : INVX0 port map( INP => n5114, ZN => n5137);
   U3826 : INVX0 port map( INP => n5114, ZN => n5138);
   U3827 : INVX0 port map( INP => n5114, ZN => n5139);
   U3828 : INVX0 port map( INP => n5114, ZN => n5140);
   U3829 : INVX0 port map( INP => n5114, ZN => n5141);
   U3830 : INVX0 port map( INP => n5115, ZN => n5142);
   U3831 : INVX0 port map( INP => n5115, ZN => n5143);
   U3832 : INVX0 port map( INP => n5115, ZN => n5144);
   U3833 : INVX0 port map( INP => n5115, ZN => n5145);
   U3834 : INVX0 port map( INP => n5115, ZN => n5146);
   U3835 : INVX0 port map( INP => n5116, ZN => n5147);
   U3836 : INVX0 port map( INP => n5116, ZN => n5148);
   U3837 : INVX0 port map( INP => n5116, ZN => n5149);
   U3838 : INVX0 port map( INP => n5116, ZN => n5150);
   U3839 : INVX0 port map( INP => n5116, ZN => n5151);
   U3840 : INVX0 port map( INP => n5493, ZN => n5528);
   U3841 : INVX0 port map( INP => n5493, ZN => n5529);
   U3842 : INVX0 port map( INP => n5451, ZN => n5486);
   U3843 : INVX0 port map( INP => n5451, ZN => n5487);
   U3844 : INVX0 port map( INP => n5159, ZN => n5194);
   U3845 : INVX0 port map( INP => n5159, ZN => n5195);
   U3846 : INVX0 port map( INP => n5117, ZN => n5152);
   U3847 : INVX0 port map( INP => n5117, ZN => n5153);
   U3848 : INVX0 port map( INP => n4988, ZN => n5007);
   U3849 : INVX0 port map( INP => n4988, ZN => n5008);
   U3850 : INVX0 port map( INP => n4988, ZN => n5009);
   U3851 : INVX0 port map( INP => n4988, ZN => n5010);
   U3852 : INVX0 port map( INP => n4988, ZN => n5011);
   U3853 : INVX0 port map( INP => n4989, ZN => n5012);
   U3854 : INVX0 port map( INP => n4989, ZN => n5013);
   U3855 : INVX0 port map( INP => n4989, ZN => n5014);
   U3856 : INVX0 port map( INP => n4989, ZN => n5015);
   U3857 : INVX0 port map( INP => n4989, ZN => n5016);
   U3858 : INVX0 port map( INP => n4990, ZN => n5017);
   U3859 : INVX0 port map( INP => n4990, ZN => n5018);
   U3860 : INVX0 port map( INP => n4990, ZN => n5019);
   U3861 : INVX0 port map( INP => n4990, ZN => n5020);
   U3862 : INVX0 port map( INP => n4990, ZN => n5021);
   U3863 : INVX0 port map( INP => n4991, ZN => n5022);
   U3864 : INVX0 port map( INP => n4991, ZN => n5023);
   U3865 : INVX0 port map( INP => n4991, ZN => n5024);
   U3866 : INVX0 port map( INP => n4991, ZN => n5025);
   U3867 : INVX0 port map( INP => n4991, ZN => n5026);
   U3868 : INVX0 port map( INP => n5072, ZN => n5091);
   U3869 : INVX0 port map( INP => n5072, ZN => n5092);
   U3870 : INVX0 port map( INP => n5072, ZN => n5093);
   U3871 : INVX0 port map( INP => n5072, ZN => n5094);
   U3872 : INVX0 port map( INP => n5073, ZN => n5095);
   U3873 : INVX0 port map( INP => n5073, ZN => n5096);
   U3874 : INVX0 port map( INP => n5073, ZN => n5097);
   U3875 : INVX0 port map( INP => n5073, ZN => n5098);
   U3876 : INVX0 port map( INP => n5073, ZN => n5099);
   U3877 : INVX0 port map( INP => n5074, ZN => n5100);
   U3878 : INVX0 port map( INP => n5074, ZN => n5101);
   U3879 : INVX0 port map( INP => n5074, ZN => n5102);
   U3880 : INVX0 port map( INP => n5074, ZN => n5103);
   U3881 : INVX0 port map( INP => n5074, ZN => n5104);
   U3882 : INVX0 port map( INP => n5075, ZN => n5105);
   U3883 : INVX0 port map( INP => n5075, ZN => n5106);
   U3884 : INVX0 port map( INP => n5075, ZN => n5107);
   U3885 : INVX0 port map( INP => n5075, ZN => n5108);
   U3886 : INVX0 port map( INP => n5075, ZN => n5109);
   U3887 : INVX0 port map( INP => n5239, ZN => n5258);
   U3888 : INVX0 port map( INP => n5239, ZN => n5259);
   U3889 : INVX0 port map( INP => n5239, ZN => n5260);
   U3890 : INVX0 port map( INP => n5239, ZN => n5261);
   U3891 : INVX0 port map( INP => n5239, ZN => n5262);
   U3892 : INVX0 port map( INP => n5240, ZN => n5263);
   U3893 : INVX0 port map( INP => n5240, ZN => n5264);
   U3894 : INVX0 port map( INP => n5240, ZN => n5265);
   U3895 : INVX0 port map( INP => n5240, ZN => n5266);
   U3896 : INVX0 port map( INP => n5240, ZN => n5267);
   U3897 : INVX0 port map( INP => n5241, ZN => n5268);
   U3898 : INVX0 port map( INP => n5241, ZN => n5269);
   U3899 : INVX0 port map( INP => n5241, ZN => n5270);
   U3900 : INVX0 port map( INP => n5241, ZN => n5271);
   U3901 : INVX0 port map( INP => n5241, ZN => n5272);
   U3902 : INVX0 port map( INP => n5242, ZN => n5273);
   U3903 : INVX0 port map( INP => n5242, ZN => n5274);
   U3904 : INVX0 port map( INP => n5242, ZN => n5275);
   U3905 : INVX0 port map( INP => n5242, ZN => n5276);
   U3906 : INVX0 port map( INP => n5242, ZN => n5277);
   U3907 : INVX0 port map( INP => n4946, ZN => n4965);
   U3908 : INVX0 port map( INP => n4946, ZN => n4966);
   U3909 : INVX0 port map( INP => n4946, ZN => n4967);
   U3910 : INVX0 port map( INP => n4946, ZN => n4968);
   U3911 : INVX0 port map( INP => n4946, ZN => n4969);
   U3912 : INVX0 port map( INP => n4947, ZN => n4970);
   U3913 : INVX0 port map( INP => n4947, ZN => n4971);
   U3914 : INVX0 port map( INP => n4947, ZN => n4972);
   U3915 : INVX0 port map( INP => n4947, ZN => n4973);
   U3916 : INVX0 port map( INP => n4947, ZN => n4974);
   U3917 : INVX0 port map( INP => n4948, ZN => n4975);
   U3918 : INVX0 port map( INP => n4948, ZN => n4976);
   U3919 : INVX0 port map( INP => n4948, ZN => n4977);
   U3920 : INVX0 port map( INP => n4948, ZN => n4978);
   U3921 : INVX0 port map( INP => n4948, ZN => n4979);
   U3922 : INVX0 port map( INP => n4949, ZN => n4980);
   U3923 : INVX0 port map( INP => n4949, ZN => n4981);
   U3924 : INVX0 port map( INP => n4949, ZN => n4982);
   U3925 : INVX0 port map( INP => n4949, ZN => n4983);
   U3926 : INVX0 port map( INP => n4949, ZN => n4984);
   U3927 : INVX0 port map( INP => n5575, ZN => n5603);
   U3928 : INVX0 port map( INP => n5575, ZN => n5604);
   U3929 : INVX0 port map( INP => n5575, ZN => n5605);
   U3930 : INVX0 port map( INP => n5573, ZN => n5592);
   U3931 : INVX0 port map( INP => n5573, ZN => n5593);
   U3932 : INVX0 port map( INP => n5573, ZN => n5594);
   U3933 : INVX0 port map( INP => n5573, ZN => n5595);
   U3934 : INVX0 port map( INP => n5573, ZN => n5596);
   U3935 : INVX0 port map( INP => n5574, ZN => n5597);
   U3936 : INVX0 port map( INP => n5574, ZN => n5598);
   U3937 : INVX0 port map( INP => n5574, ZN => n5599);
   U3938 : INVX0 port map( INP => n5574, ZN => n5601);
   U3939 : INVX0 port map( INP => n5575, ZN => n5602);
   U3940 : INVX0 port map( INP => n5575, ZN => n5606);
   U3941 : INVX0 port map( INP => n5576, ZN => n5607);
   U3942 : INVX0 port map( INP => n5576, ZN => n5608);
   U3943 : INVX0 port map( INP => n5576, ZN => n5609);
   U3944 : INVX0 port map( INP => n5576, ZN => n5610);
   U3945 : INVX0 port map( INP => n5576, ZN => n5611);
   U3946 : INVX0 port map( INP => n5577, ZN => n5612);
   U3947 : INVX0 port map( INP => n5577, ZN => n5613);
   U3948 : INVX0 port map( INP => n5327, ZN => n5364);
   U3949 : INVX0 port map( INP => n5410, ZN => n5446);
   U3950 : INVX0 port map( INP => n5493, ZN => n5530);
   U3951 : INVX0 port map( INP => n5451, ZN => n5488);
   U3952 : INVX0 port map( INP => n5159, ZN => n5196);
   U3953 : INVX0 port map( INP => n5117, ZN => n5154);
   U3954 : INVX0 port map( INP => n5577, ZN => n5614);
   U3955 : INVX0 port map( INP => n5536, ZN => n5532);
   U3956 : INVX0 port map( INP => n5536, ZN => n5533);
   U3957 : INVX0 port map( INP => n5536, ZN => n5531);
   U3958 : INVX0 port map( INP => n5536, ZN => n5534);
   U3959 : INVX0 port map( INP => n5370, ZN => n5365);
   U3960 : INVX0 port map( INP => n5370, ZN => n5366);
   U3961 : INVX0 port map( INP => n5370, ZN => n5367);
   U3962 : INVX0 port map( INP => n5370, ZN => n5368);
   U3963 : INVX0 port map( INP => n4992, ZN => n5027);
   U3964 : INVX0 port map( INP => n4992, ZN => n5028);
   U3965 : INVX0 port map( INP => n5076, ZN => n5110);
   U3966 : INVX0 port map( INP => n5076, ZN => n5111);
   U3967 : INVX0 port map( INP => n5243, ZN => n5278);
   U3968 : INVX0 port map( INP => n5243, ZN => n5279);
   U3969 : INVX0 port map( INP => n4950, ZN => n4985);
   U3970 : INVX0 port map( INP => n4950, ZN => n4986);
   U3971 : INVX0 port map( INP => n5281, ZN => n5300);
   U3972 : INVX0 port map( INP => n5281, ZN => n5301);
   U3973 : INVX0 port map( INP => n5281, ZN => n5302);
   U3974 : INVX0 port map( INP => n5281, ZN => n5303);
   U3975 : INVX0 port map( INP => n5281, ZN => n5304);
   U3976 : INVX0 port map( INP => n5282, ZN => n5305);
   U3977 : INVX0 port map( INP => n5282, ZN => n5306);
   U3978 : INVX0 port map( INP => n5282, ZN => n5307);
   U3979 : INVX0 port map( INP => n5282, ZN => n5308);
   U3980 : INVX0 port map( INP => n5282, ZN => n5309);
   U3981 : INVX0 port map( INP => n5283, ZN => n5310);
   U3982 : INVX0 port map( INP => n5283, ZN => n5311);
   U3983 : INVX0 port map( INP => n5283, ZN => n5312);
   U3984 : INVX0 port map( INP => n5283, ZN => n5313);
   U3985 : INVX0 port map( INP => n5283, ZN => n5314);
   U3986 : INVX0 port map( INP => n5284, ZN => n5315);
   U3987 : INVX0 port map( INP => n5284, ZN => n5316);
   U3988 : INVX0 port map( INP => n5284, ZN => n5317);
   U3989 : INVX0 port map( INP => n5284, ZN => n5318);
   U3990 : INVX0 port map( INP => n5284, ZN => n5319);
   U3991 : INVX0 port map( INP => n5285, ZN => n5320);
   U3992 : INVX0 port map( INP => n5285, ZN => n5321);
   U3993 : INVX0 port map( INP => n4992, ZN => n5029);
   U3994 : INVX0 port map( INP => n5076, ZN => n5112);
   U3995 : INVX0 port map( INP => n5243, ZN => n5280);
   U3996 : INVX0 port map( INP => n4950, ZN => n4987);
   U3997 : INVX0 port map( INP => n5285, ZN => n5322);
   U3998 : INVX0 port map( INP => n5035, ZN => n5034);
   U3999 : INVX0 port map( INP => n5202, ZN => n5201);
   U4000 : INVX0 port map( INP => n5536, ZN => n5535);
   U4001 : INVX0 port map( INP => n5370, ZN => n5369);
   U4002 : INVX0 port map( INP => n26, ZN => n5507);
   U4003 : INVX0 port map( INP => n28, ZN => n5465);
   U4004 : INVX0 port map( INP => n40, ZN => n5173);
   U4005 : INVX0 port map( INP => n41, ZN => n5131);
   U4006 : INVX0 port map( INP => n21, ZN => n5590);
   U4007 : INVX0 port map( INP => n44, ZN => n5006);
   U4008 : INVX0 port map( INP => n42, ZN => n5090);
   U4009 : INVX0 port map( INP => n36, ZN => n5257);
   U4010 : INVX0 port map( INP => n46, ZN => n4964);
   U4011 : INVX0 port map( INP => n26, ZN => n5506);
   U4012 : INVX0 port map( INP => n28, ZN => n5464);
   U4013 : INVX0 port map( INP => n40, ZN => n5172);
   U4014 : INVX0 port map( INP => n41, ZN => n5130);
   U4015 : INVX0 port map( INP => n44, ZN => n5005);
   U4016 : INVX0 port map( INP => n42, ZN => n5089);
   U4017 : INVX0 port map( INP => n36, ZN => n5256);
   U4018 : INVX0 port map( INP => n46, ZN => n4963);
   U4019 : INVX0 port map( INP => n21, ZN => n5591);
   U4020 : INVX0 port map( INP => n32, ZN => n5340);
   U4021 : INVX0 port map( INP => n29, ZN => n5423);
   U4022 : INVX0 port map( INP => n35, ZN => n5299);
   U4023 : INVX0 port map( INP => n35, ZN => n5298);
   U4024 : INVX0 port map( INP => n5578, ZN => n5574);
   U4025 : INVX0 port map( INP => n5578, ZN => n5575);
   U4026 : INVX0 port map( INP => n5578, ZN => n5573);
   U4027 : INVX0 port map( INP => n5578, ZN => n5576);
   U4028 : INVX0 port map( INP => n5328, ZN => n5323);
   U4029 : INVX0 port map( INP => n5328, ZN => n5324);
   U4030 : INVX0 port map( INP => n5328, ZN => n5325);
   U4031 : INVX0 port map( INP => n5328, ZN => n5326);
   U4032 : INVX0 port map( INP => n5411, ZN => n5406);
   U4033 : INVX0 port map( INP => n5411, ZN => n5407);
   U4034 : INVX0 port map( INP => n5411, ZN => n5408);
   U4035 : INVX0 port map( INP => n5411, ZN => n5409);
   U4036 : INVX0 port map( INP => n5494, ZN => n5489);
   U4037 : INVX0 port map( INP => n5494, ZN => n5490);
   U4038 : INVX0 port map( INP => n5494, ZN => n5491);
   U4039 : INVX0 port map( INP => n5494, ZN => n5492);
   U4040 : INVX0 port map( INP => n5452, ZN => n5447);
   U4041 : INVX0 port map( INP => n5452, ZN => n5448);
   U4042 : INVX0 port map( INP => n5452, ZN => n5449);
   U4043 : INVX0 port map( INP => n5452, ZN => n5450);
   U4044 : INVX0 port map( INP => n5160, ZN => n5155);
   U4045 : INVX0 port map( INP => n5160, ZN => n5156);
   U4046 : INVX0 port map( INP => n5160, ZN => n5157);
   U4047 : INVX0 port map( INP => n5160, ZN => n5158);
   U4048 : INVX0 port map( INP => n5118, ZN => n5113);
   U4049 : INVX0 port map( INP => n5118, ZN => n5114);
   U4050 : INVX0 port map( INP => n5118, ZN => n5115);
   U4051 : INVX0 port map( INP => n5118, ZN => n5116);
   U4052 : INVX0 port map( INP => n4993, ZN => n4988);
   U4053 : INVX0 port map( INP => n4993, ZN => n4989);
   U4054 : INVX0 port map( INP => n4993, ZN => n4990);
   U4055 : INVX0 port map( INP => n4993, ZN => n4991);
   U4056 : INVX0 port map( INP => n5077, ZN => n5072);
   U4057 : INVX0 port map( INP => n5077, ZN => n5073);
   U4058 : INVX0 port map( INP => n5077, ZN => n5074);
   U4059 : INVX0 port map( INP => n5077, ZN => n5075);
   U4060 : INVX0 port map( INP => n5244, ZN => n5239);
   U4061 : INVX0 port map( INP => n5244, ZN => n5240);
   U4062 : INVX0 port map( INP => n5244, ZN => n5241);
   U4063 : INVX0 port map( INP => n5244, ZN => n5242);
   U4064 : INVX0 port map( INP => n4951, ZN => n4946);
   U4065 : INVX0 port map( INP => n4951, ZN => n4947);
   U4066 : INVX0 port map( INP => n4951, ZN => n4948);
   U4067 : INVX0 port map( INP => n4951, ZN => n4949);
   U4068 : INVX0 port map( INP => n38, ZN => n5202);
   U4069 : INVX0 port map( INP => n43, ZN => n5035);
   U4070 : INVX0 port map( INP => n5578, ZN => n5577);
   U4071 : INVX0 port map( INP => n5328, ZN => n5327);
   U4072 : INVX0 port map( INP => n5411, ZN => n5410);
   U4073 : INVX0 port map( INP => n5494, ZN => n5493);
   U4074 : INVX0 port map( INP => n5452, ZN => n5451);
   U4075 : INVX0 port map( INP => n5160, ZN => n5159);
   U4076 : INVX0 port map( INP => n5118, ZN => n5117);
   U4077 : INVX0 port map( INP => n5286, ZN => n5281);
   U4078 : INVX0 port map( INP => n5286, ZN => n5282);
   U4079 : INVX0 port map( INP => n5286, ZN => n5283);
   U4080 : INVX0 port map( INP => n5286, ZN => n5284);
   U4081 : INVX0 port map( INP => n31, ZN => n5370);
   U4082 : INVX0 port map( INP => n24, ZN => n5536);
   U4083 : INVX0 port map( INP => n4993, ZN => n4992);
   U4084 : INVX0 port map( INP => n5077, ZN => n5076);
   U4085 : INVX0 port map( INP => n5244, ZN => n5243);
   U4086 : INVX0 port map( INP => n4951, ZN => n4950);
   U4087 : INVX0 port map( INP => n5286, ZN => n5285);
   U4088 : NBUFFX2 port map( INP => n4743, Z => n4929);
   U4089 : NBUFFX2 port map( INP => n4743, Z => n4928);
   U4090 : NBUFFX2 port map( INP => n4744, Z => n4932);
   U4091 : NBUFFX2 port map( INP => n4744, Z => n4931);
   U4092 : NBUFFX2 port map( INP => n4743, Z => n4930);
   U4093 : NBUFFX2 port map( INP => n4745, Z => n4936);
   U4094 : NBUFFX2 port map( INP => n4745, Z => n4935);
   U4095 : NBUFFX2 port map( INP => n4745, Z => n4934);
   U4096 : NBUFFX2 port map( INP => n4744, Z => n4933);
   U4097 : NBUFFX2 port map( INP => n4740, Z => n4920);
   U4098 : NBUFFX2 port map( INP => n4740, Z => n4919);
   U4099 : NBUFFX2 port map( INP => n4741, Z => n4923);
   U4100 : NBUFFX2 port map( INP => n4741, Z => n4922);
   U4101 : NBUFFX2 port map( INP => n4740, Z => n4921);
   U4102 : NBUFFX2 port map( INP => n4742, Z => n4927);
   U4103 : NBUFFX2 port map( INP => n4742, Z => n4926);
   U4104 : NBUFFX2 port map( INP => n4742, Z => n4925);
   U4105 : NBUFFX2 port map( INP => n4741, Z => n4924);
   U4106 : NBUFFX2 port map( INP => n4737, Z => n4911);
   U4107 : NBUFFX2 port map( INP => n4737, Z => n4910);
   U4108 : NBUFFX2 port map( INP => n4738, Z => n4914);
   U4109 : NBUFFX2 port map( INP => n4738, Z => n4913);
   U4110 : NBUFFX2 port map( INP => n4737, Z => n4912);
   U4111 : NBUFFX2 port map( INP => n4739, Z => n4918);
   U4112 : NBUFFX2 port map( INP => n4739, Z => n4917);
   U4113 : NBUFFX2 port map( INP => n4739, Z => n4916);
   U4114 : NBUFFX2 port map( INP => n4738, Z => n4915);
   U4115 : NBUFFX2 port map( INP => n4734, Z => n4902);
   U4116 : NBUFFX2 port map( INP => n4734, Z => n4901);
   U4117 : NBUFFX2 port map( INP => n4735, Z => n4905);
   U4118 : NBUFFX2 port map( INP => n4735, Z => n4904);
   U4119 : NBUFFX2 port map( INP => n4734, Z => n4903);
   U4120 : NBUFFX2 port map( INP => n4736, Z => n4909);
   U4121 : NBUFFX2 port map( INP => n4736, Z => n4908);
   U4122 : NBUFFX2 port map( INP => n4736, Z => n4907);
   U4123 : NBUFFX2 port map( INP => n4735, Z => n4906);
   U4124 : NBUFFX2 port map( INP => n4731, Z => n4893);
   U4125 : NBUFFX2 port map( INP => n4731, Z => n4892);
   U4126 : NBUFFX2 port map( INP => n4732, Z => n4896);
   U4127 : NBUFFX2 port map( INP => n4732, Z => n4895);
   U4128 : NBUFFX2 port map( INP => n4731, Z => n4894);
   U4129 : NBUFFX2 port map( INP => n4733, Z => n4900);
   U4130 : NBUFFX2 port map( INP => n4733, Z => n4899);
   U4131 : NBUFFX2 port map( INP => n4733, Z => n4898);
   U4132 : NBUFFX2 port map( INP => n4732, Z => n4897);
   U4133 : NBUFFX2 port map( INP => n4728, Z => n4884);
   U4134 : NBUFFX2 port map( INP => n4728, Z => n4883);
   U4135 : NBUFFX2 port map( INP => n4729, Z => n4887);
   U4136 : NBUFFX2 port map( INP => n4729, Z => n4886);
   U4137 : NBUFFX2 port map( INP => n4728, Z => n4885);
   U4138 : NBUFFX2 port map( INP => n4730, Z => n4891);
   U4139 : NBUFFX2 port map( INP => n4730, Z => n4890);
   U4140 : NBUFFX2 port map( INP => n4730, Z => n4889);
   U4141 : NBUFFX2 port map( INP => n4729, Z => n4888);
   U4142 : NBUFFX2 port map( INP => n4725, Z => n4875);
   U4143 : NBUFFX2 port map( INP => n4725, Z => n4874);
   U4144 : NBUFFX2 port map( INP => n4726, Z => n4878);
   U4145 : NBUFFX2 port map( INP => n4726, Z => n4877);
   U4146 : NBUFFX2 port map( INP => n4725, Z => n4876);
   U4147 : NBUFFX2 port map( INP => n4727, Z => n4882);
   U4148 : NBUFFX2 port map( INP => n4727, Z => n4881);
   U4149 : NBUFFX2 port map( INP => n4727, Z => n4880);
   U4150 : NBUFFX2 port map( INP => n4726, Z => n4879);
   U4151 : NBUFFX2 port map( INP => n4722, Z => n4866);
   U4152 : NBUFFX2 port map( INP => n4722, Z => n4865);
   U4153 : NBUFFX2 port map( INP => n4723, Z => n4869);
   U4154 : NBUFFX2 port map( INP => n4723, Z => n4868);
   U4155 : NBUFFX2 port map( INP => n4722, Z => n4867);
   U4156 : NBUFFX2 port map( INP => n4724, Z => n4873);
   U4157 : NBUFFX2 port map( INP => n4724, Z => n4872);
   U4158 : NBUFFX2 port map( INP => n4724, Z => n4871);
   U4159 : NBUFFX2 port map( INP => n4723, Z => n4870);
   U4160 : NBUFFX2 port map( INP => n4719, Z => n4857);
   U4161 : NBUFFX2 port map( INP => n4719, Z => n4856);
   U4162 : NBUFFX2 port map( INP => n4720, Z => n4860);
   U4163 : NBUFFX2 port map( INP => n4720, Z => n4859);
   U4164 : NBUFFX2 port map( INP => n4719, Z => n4858);
   U4165 : NBUFFX2 port map( INP => n4721, Z => n4864);
   U4166 : NBUFFX2 port map( INP => n4721, Z => n4863);
   U4167 : NBUFFX2 port map( INP => n4721, Z => n4862);
   U4168 : NBUFFX2 port map( INP => n4720, Z => n4861);
   U4169 : NBUFFX2 port map( INP => n4716, Z => n4848);
   U4170 : NBUFFX2 port map( INP => n4716, Z => n4847);
   U4171 : NBUFFX2 port map( INP => n4717, Z => n4851);
   U4172 : NBUFFX2 port map( INP => n4717, Z => n4850);
   U4173 : NBUFFX2 port map( INP => n4716, Z => n4849);
   U4174 : NBUFFX2 port map( INP => n4718, Z => n4855);
   U4175 : NBUFFX2 port map( INP => n4718, Z => n4854);
   U4176 : NBUFFX2 port map( INP => n4718, Z => n4853);
   U4177 : NBUFFX2 port map( INP => n4717, Z => n4852);
   U4178 : NBUFFX2 port map( INP => n4713, Z => n4839);
   U4179 : NBUFFX2 port map( INP => n4713, Z => n4838);
   U4180 : NBUFFX2 port map( INP => n4714, Z => n4842);
   U4181 : NBUFFX2 port map( INP => n4714, Z => n4841);
   U4182 : NBUFFX2 port map( INP => n4713, Z => n4840);
   U4183 : NBUFFX2 port map( INP => n4715, Z => n4846);
   U4184 : NBUFFX2 port map( INP => n4715, Z => n4845);
   U4185 : NBUFFX2 port map( INP => n4715, Z => n4844);
   U4186 : NBUFFX2 port map( INP => n4714, Z => n4843);
   U4187 : NBUFFX2 port map( INP => n4710, Z => n4830);
   U4188 : NBUFFX2 port map( INP => n4710, Z => n4829);
   U4189 : NBUFFX2 port map( INP => n4711, Z => n4833);
   U4190 : NBUFFX2 port map( INP => n4711, Z => n4832);
   U4191 : NBUFFX2 port map( INP => n4710, Z => n4831);
   U4192 : NBUFFX2 port map( INP => n4712, Z => n4837);
   U4193 : NBUFFX2 port map( INP => n4712, Z => n4836);
   U4194 : NBUFFX2 port map( INP => n4712, Z => n4835);
   U4195 : NBUFFX2 port map( INP => n4711, Z => n4834);
   U4196 : NBUFFX2 port map( INP => n4707, Z => n4821);
   U4197 : NBUFFX2 port map( INP => n4707, Z => n4820);
   U4198 : NBUFFX2 port map( INP => n4708, Z => n4824);
   U4199 : NBUFFX2 port map( INP => n4708, Z => n4823);
   U4200 : NBUFFX2 port map( INP => n4707, Z => n4822);
   U4201 : NBUFFX2 port map( INP => n4709, Z => n4828);
   U4202 : NBUFFX2 port map( INP => n4709, Z => n4827);
   U4203 : NBUFFX2 port map( INP => n4709, Z => n4826);
   U4204 : NBUFFX2 port map( INP => n4708, Z => n4825);
   U4205 : NBUFFX2 port map( INP => n4704, Z => n4812);
   U4206 : NBUFFX2 port map( INP => n4704, Z => n4811);
   U4207 : NBUFFX2 port map( INP => n4705, Z => n4815);
   U4208 : NBUFFX2 port map( INP => n4705, Z => n4814);
   U4209 : NBUFFX2 port map( INP => n4704, Z => n4813);
   U4210 : NBUFFX2 port map( INP => n4706, Z => n4819);
   U4211 : NBUFFX2 port map( INP => n4706, Z => n4818);
   U4212 : NBUFFX2 port map( INP => n4706, Z => n4817);
   U4213 : NBUFFX2 port map( INP => n4705, Z => n4816);
   U4214 : NBUFFX2 port map( INP => n4701, Z => n4803);
   U4215 : NBUFFX2 port map( INP => n4701, Z => n4802);
   U4216 : NBUFFX2 port map( INP => n4702, Z => n4806);
   U4217 : NBUFFX2 port map( INP => n4702, Z => n4805);
   U4218 : NBUFFX2 port map( INP => n4701, Z => n4804);
   U4219 : NBUFFX2 port map( INP => n4703, Z => n4810);
   U4220 : NBUFFX2 port map( INP => n4703, Z => n4809);
   U4221 : NBUFFX2 port map( INP => n4703, Z => n4808);
   U4222 : NBUFFX2 port map( INP => n4702, Z => n4807);
   U4223 : NBUFFX2 port map( INP => n4698, Z => n4794);
   U4224 : NBUFFX2 port map( INP => n4698, Z => n4793);
   U4225 : NBUFFX2 port map( INP => n4699, Z => n4797);
   U4226 : NBUFFX2 port map( INP => n4699, Z => n4796);
   U4227 : NBUFFX2 port map( INP => n4698, Z => n4795);
   U4228 : NBUFFX2 port map( INP => n4700, Z => n4801);
   U4229 : NBUFFX2 port map( INP => n4700, Z => n4800);
   U4230 : NBUFFX2 port map( INP => n4700, Z => n4799);
   U4231 : NBUFFX2 port map( INP => n4699, Z => n4798);
   U4232 : NBUFFX2 port map( INP => n4695, Z => n4785);
   U4233 : NBUFFX2 port map( INP => n4695, Z => n4784);
   U4234 : NBUFFX2 port map( INP => n4696, Z => n4788);
   U4235 : NBUFFX2 port map( INP => n4696, Z => n4787);
   U4236 : NBUFFX2 port map( INP => n4695, Z => n4786);
   U4237 : NBUFFX2 port map( INP => n4697, Z => n4792);
   U4238 : NBUFFX2 port map( INP => n4697, Z => n4791);
   U4239 : NBUFFX2 port map( INP => n4697, Z => n4790);
   U4240 : NBUFFX2 port map( INP => n4696, Z => n4789);
   U4241 : NBUFFX2 port map( INP => n4692, Z => n4777);
   U4242 : NBUFFX2 port map( INP => n4692, Z => n4776);
   U4243 : NBUFFX2 port map( INP => n4692, Z => n4775);
   U4244 : NBUFFX2 port map( INP => n4693, Z => n4780);
   U4245 : NBUFFX2 port map( INP => n4693, Z => n4779);
   U4246 : NBUFFX2 port map( INP => n4693, Z => n4778);
   U4247 : NBUFFX2 port map( INP => n4694, Z => n4783);
   U4248 : NBUFFX2 port map( INP => n4694, Z => n4782);
   U4249 : NBUFFX2 port map( INP => n4694, Z => n4781);
   U4250 : INVX0 port map( INP => n3340, ZN => n3464);
   U4251 : NBUFFX2 port map( INP => n3344, Z => n3444);
   U4252 : NBUFFX2 port map( INP => n3344, Z => n3442);
   U4253 : NBUFFX2 port map( INP => n3344, Z => n3445);
   U4254 : DELLN1X2 port map( INP => n3346, Z => n3376);
   U4255 : DELLN1X2 port map( INP => n3342, Z => n3367);
   U4256 : DELLN1X2 port map( INP => n3346, Z => n3378);
   U4257 : DELLN1X2 port map( INP => n3342, Z => n3368);
   U4258 : DELLN1X2 port map( INP => n3342, Z => n3365);
   U4259 : DELLN1X2 port map( INP => n3346, Z => n3379);
   U4260 : DELLN1X2 port map( INP => n3342, Z => n3366);
   U4261 : DELLN1X2 port map( INP => n3342, Z => n3361);
   U4262 : DELLN1X2 port map( INP => n3342, Z => n3369);
   U4263 : DELLN1X2 port map( INP => n3356, Z => n3396);
   U4264 : DELLN1X2 port map( INP => n3356, Z => n3398);
   U4265 : DELLN1X2 port map( INP => n3356, Z => n3392);
   U4266 : DELLN1X2 port map( INP => n3356, Z => n3397);
   U4267 : DELLN1X2 port map( INP => n3356, Z => n3400);
   U4268 : DELLN1X2 port map( INP => n3351, Z => n3388);
   U4269 : DELLN1X2 port map( INP => n3351, Z => n3387);
   U4270 : DELLN1X2 port map( INP => n3351, Z => n3384);
   U4271 : DELLN1X2 port map( INP => n3351, Z => n3386);
   U4272 : DELLN1X2 port map( INP => n3342, Z => n3362);
   U4273 : DELLN1X2 port map( INP => n3342, Z => n3370);
   U4274 : DELLN1X2 port map( INP => n3346, Z => n3381);
   U4275 : NBUFFX2 port map( INP => n3427, Z => n3425);
   U4276 : NBUFFX2 port map( INP => n3427, Z => n3421);
   U4277 : NBUFFX2 port map( INP => n3427, Z => n3426);
   U4278 : NBUFFX2 port map( INP => n3427, Z => n3422);
   U4279 : NBUFFX2 port map( INP => n3427, Z => n3424);
   U4280 : DELLN1X2 port map( INP => n4494, Z => n4562);
   U4281 : NBUFFX2 port map( INP => n4494, Z => n4568);
   U4282 : NBUFFX2 port map( INP => n4494, Z => n4569);
   U4283 : NBUFFX2 port map( INP => n4494, Z => n4565);
   U4284 : NBUFFX2 port map( INP => n4494, Z => n4567);
   U4285 : NBUFFX2 port map( INP => n4494, Z => n4564);
   U4286 : NBUFFX2 port map( INP => n4494, Z => n4563);
   U4287 : NBUFFX2 port map( INP => n4504, Z => n4653);
   U4288 : NBUFFX2 port map( INP => n4495, Z => n4576);
   U4289 : DELLN1X2 port map( INP => n4507, Z => n4672);
   U4290 : DELLN1X2 port map( INP => n4502, Z => n4628);
   U4291 : DELLN1X2 port map( INP => n4492, Z => n4540);
   U4292 : DELLN1X2 port map( INP => n4507, Z => n4676);
   U4293 : DELLN1X2 port map( INP => n4502, Z => n4632);
   U4294 : DELLN1X2 port map( INP => n4492, Z => n4544);
   U4295 : DELLN1X2 port map( INP => n4497, Z => n4584);
   U4296 : DELLN1X2 port map( INP => n4497, Z => n4588);
   U4297 : DELLN1X2 port map( INP => n4507, Z => n4671);
   U4298 : DELLN1X2 port map( INP => n4507, Z => n4680);
   U4299 : DELLN1X2 port map( INP => n4502, Z => n4627);
   U4300 : DELLN1X2 port map( INP => n4492, Z => n4539);
   U4301 : DELLN1X2 port map( INP => n4502, Z => n4636);
   U4302 : DELLN1X2 port map( INP => n4492, Z => n4548);
   U4303 : NBUFFX2 port map( INP => n4507, Z => n4677);
   U4304 : NBUFFX2 port map( INP => n4507, Z => n4674);
   U4305 : NBUFFX2 port map( INP => n4507, Z => n4675);
   U4306 : NBUFFX2 port map( INP => n4507, Z => n4673);
   U4307 : NBUFFX2 port map( INP => n4502, Z => n4633);
   U4308 : NBUFFX2 port map( INP => n4502, Z => n4630);
   U4309 : NBUFFX2 port map( INP => n4502, Z => n4631);
   U4310 : NBUFFX2 port map( INP => n4502, Z => n4629);
   U4311 : NBUFFX2 port map( INP => n4492, Z => n4545);
   U4312 : NBUFFX2 port map( INP => n4492, Z => n4542);
   U4313 : NBUFFX2 port map( INP => n4492, Z => n4543);
   U4314 : NBUFFX2 port map( INP => n4492, Z => n4541);
   U4315 : NBUFFX2 port map( INP => n4497, Z => n4590);
   U4316 : NBUFFX2 port map( INP => n4497, Z => n4591);
   U4317 : NBUFFX2 port map( INP => n4497, Z => n4587);
   U4318 : NBUFFX2 port map( INP => n4497, Z => n4589);
   U4319 : NBUFFX2 port map( INP => n4497, Z => n4586);
   U4320 : NBUFFX2 port map( INP => n4497, Z => n4585);
   U4321 : DELLN1X2 port map( INP => n4494, Z => n4566);
   U4322 : DELLN1X2 port map( INP => n4499, Z => n4606);
   U4323 : DELLN1X2 port map( INP => n4504, Z => n4650);
   U4324 : DELLN1X2 port map( INP => n4489, Z => n4518);
   U4325 : DELLN1X2 port map( INP => n4499, Z => n4610);
   U4326 : DELLN1X2 port map( INP => n4504, Z => n4654);
   U4327 : DELLN1X2 port map( INP => n4489, Z => n4522);
   U4328 : NBUFFX2 port map( INP => n4504, Z => n4655);
   U4329 : NBUFFX2 port map( INP => n4504, Z => n4652);
   U4330 : NBUFFX2 port map( INP => n4504, Z => n4651);
   U4331 : NBUFFX2 port map( INP => n4499, Z => n4609);
   U4332 : NBUFFX2 port map( INP => n4489, Z => n4521);
   U4333 : NBUFFX2 port map( INP => n4499, Z => n4611);
   U4334 : NBUFFX2 port map( INP => n4499, Z => n4608);
   U4335 : NBUFFX2 port map( INP => n4499, Z => n4607);
   U4336 : NBUFFX2 port map( INP => n4489, Z => n4523);
   U4337 : NBUFFX2 port map( INP => n4489, Z => n4520);
   U4338 : NBUFFX2 port map( INP => n4489, Z => n4519);
   U4339 : DELLN1X2 port map( INP => n4508, Z => n4683);
   U4340 : DELLN1X2 port map( INP => n4508, Z => n4687);
   U4341 : DELLN1X2 port map( INP => n4498, Z => n4595);
   U4342 : DELLN1X2 port map( INP => n4498, Z => n4599);
   U4343 : NBUFFX2 port map( INP => n4508, Z => n4688);
   U4344 : NBUFFX2 port map( INP => n4508, Z => n4685);
   U4345 : NBUFFX2 port map( INP => n4508, Z => n4686);
   U4346 : NBUFFX2 port map( INP => n4508, Z => n4684);
   U4347 : NBUFFX2 port map( INP => n4498, Z => n4601);
   U4348 : NBUFFX2 port map( INP => n4498, Z => n4602);
   U4349 : NBUFFX2 port map( INP => n4493, Z => n4554);
   U4350 : NBUFFX2 port map( INP => n4498, Z => n4598);
   U4351 : NBUFFX2 port map( INP => n4498, Z => n4600);
   U4352 : NBUFFX2 port map( INP => n4498, Z => n4597);
   U4353 : NBUFFX2 port map( INP => n4498, Z => n4596);
   U4354 : DELLN1X2 port map( INP => n4505, Z => n4661);
   U4355 : DELLN1X2 port map( INP => n4490, Z => n4529);
   U4356 : DELLN1X2 port map( INP => n4505, Z => n4665);
   U4357 : DELLN1X2 port map( INP => n4490, Z => n4533);
   U4358 : DELLN1X2 port map( INP => n4495, Z => n4573);
   U4359 : DELLN1X2 port map( INP => n4495, Z => n4577);
   U4360 : NBUFFX2 port map( INP => n4495, Z => n4579);
   U4361 : NBUFFX2 port map( INP => n4495, Z => n4580);
   U4362 : NBUFFX2 port map( INP => n4505, Z => n4664);
   U4363 : NBUFFX2 port map( INP => n4495, Z => n4578);
   U4364 : NBUFFX2 port map( INP => n4495, Z => n4575);
   U4365 : NBUFFX2 port map( INP => n4495, Z => n4574);
   U4366 : NBUFFX2 port map( INP => n4505, Z => n4666);
   U4367 : NBUFFX2 port map( INP => n4505, Z => n4663);
   U4368 : NBUFFX2 port map( INP => n4505, Z => n4662);
   U4369 : NBUFFX2 port map( INP => n4490, Z => n4532);
   U4370 : NBUFFX2 port map( INP => n4490, Z => n4534);
   U4371 : NBUFFX2 port map( INP => n4490, Z => n4531);
   U4372 : NBUFFX2 port map( INP => n4490, Z => n4530);
   U4373 : NBUFFX2 port map( INP => n4500, Z => n4620);
   U4374 : NBUFFX2 port map( INP => n4494, Z => n4560);
   U4375 : NBUFFX2 port map( INP => n4504, Z => n4648);
   U4376 : NBUFFX2 port map( INP => n4499, Z => n4604);
   U4377 : NBUFFX2 port map( INP => n4489, Z => n4516);
   U4378 : NBUFFX2 port map( INP => n4495, Z => n4571);
   U4379 : NBUFFX2 port map( INP => n4505, Z => n4659);
   U4380 : NBUFFX2 port map( INP => n4490, Z => n4527);
   U4381 : DELLN1X2 port map( INP => n4493, Z => n4551);
   U4382 : DELLN1X2 port map( INP => n4503, Z => n4639);
   U4383 : DELLN1X2 port map( INP => n4493, Z => n4555);
   U4384 : DELLN1X2 port map( INP => n4503, Z => n4643);
   U4385 : DELLN1X2 port map( INP => n4493, Z => n4550);
   U4386 : DELLN1X2 port map( INP => n4493, Z => n4559);
   U4387 : DELLN1X2 port map( INP => n4503, Z => n4638);
   U4388 : DELLN1X2 port map( INP => n4503, Z => n4647);
   U4389 : NBUFFX2 port map( INP => n4493, Z => n4556);
   U4390 : NBUFFX2 port map( INP => n4493, Z => n4553);
   U4391 : NBUFFX2 port map( INP => n4493, Z => n4552);
   U4392 : NBUFFX2 port map( INP => n4503, Z => n4642);
   U4393 : NBUFFX2 port map( INP => n4503, Z => n4644);
   U4394 : NBUFFX2 port map( INP => n4503, Z => n4641);
   U4395 : NBUFFX2 port map( INP => n4503, Z => n4640);
   U4396 : DELLN1X2 port map( INP => n4500, Z => n4617);
   U4397 : DELLN1X2 port map( INP => n4500, Z => n4621);
   U4398 : NBUFFX2 port map( INP => n4500, Z => n4622);
   U4399 : NBUFFX2 port map( INP => n4500, Z => n4619);
   U4400 : NBUFFX2 port map( INP => n4500, Z => n4618);
   U4401 : NBUFFX2 port map( INP => n4507, Z => n4670);
   U4402 : NBUFFX2 port map( INP => n4502, Z => n4626);
   U4403 : NBUFFX2 port map( INP => n4492, Z => n4538);
   U4404 : NBUFFX2 port map( INP => n4497, Z => n4582);
   U4405 : NBUFFX2 port map( INP => n4508, Z => n4681);
   U4406 : NBUFFX2 port map( INP => n4493, Z => n4549);
   U4407 : NBUFFX2 port map( INP => n4498, Z => n4593);
   U4408 : NBUFFX2 port map( INP => n4500, Z => n4615);
   U4409 : NBUFFX2 port map( INP => n4503, Z => n4637);
   U4410 : INVX0 port map( INP => n21, ZN => n5578);
   U4411 : INVX0 port map( INP => n32, ZN => n5328);
   U4412 : INVX0 port map( INP => n29, ZN => n5411);
   U4413 : INVX0 port map( INP => n28, ZN => n5452);
   U4414 : INVX0 port map( INP => n26, ZN => n5494);
   U4415 : INVX0 port map( INP => n40, ZN => n5160);
   U4416 : INVX0 port map( INP => n41, ZN => n5118);
   U4417 : INVX0 port map( INP => n36, ZN => n5244);
   U4418 : INVX0 port map( INP => n44, ZN => n4993);
   U4419 : INVX0 port map( INP => n42, ZN => n5077);
   U4420 : INVX0 port map( INP => n46, ZN => n4951);
   U4421 : INVX0 port map( INP => n35, ZN => n5286);
   U4422 : NBUFFX2 port map( INP => n4746, Z => n4938);
   U4423 : NBUFFX2 port map( INP => n4746, Z => n4937);
   U4424 : NBUFFX2 port map( INP => n4747, Z => n4941);
   U4425 : NBUFFX2 port map( INP => n4747, Z => n4940);
   U4426 : NBUFFX2 port map( INP => n4746, Z => n4939);
   U4427 : NBUFFX2 port map( INP => n4748, Z => n4944);
   U4428 : NBUFFX2 port map( INP => n4748, Z => n4943);
   U4429 : NBUFFX2 port map( INP => n4747, Z => n4942);
   U4430 : NBUFFX2 port map( INP => n4748, Z => n4945);
   U4431 : NBUFFX2 port map( INP => n4750, Z => n4743);
   U4432 : NBUFFX2 port map( INP => n4750, Z => n4745);
   U4433 : NBUFFX2 port map( INP => n4750, Z => n4744);
   U4434 : NBUFFX2 port map( INP => n4751, Z => n4740);
   U4435 : NBUFFX2 port map( INP => n4751, Z => n4742);
   U4436 : NBUFFX2 port map( INP => n4751, Z => n4741);
   U4437 : NBUFFX2 port map( INP => n4752, Z => n4737);
   U4438 : NBUFFX2 port map( INP => n4752, Z => n4739);
   U4439 : NBUFFX2 port map( INP => n4752, Z => n4738);
   U4440 : NBUFFX2 port map( INP => n4753, Z => n4734);
   U4441 : NBUFFX2 port map( INP => n4753, Z => n4736);
   U4442 : NBUFFX2 port map( INP => n4753, Z => n4735);
   U4443 : NBUFFX2 port map( INP => n4754, Z => n4731);
   U4444 : NBUFFX2 port map( INP => n4754, Z => n4733);
   U4445 : NBUFFX2 port map( INP => n4754, Z => n4732);
   U4446 : NBUFFX2 port map( INP => n4755, Z => n4728);
   U4447 : NBUFFX2 port map( INP => n4755, Z => n4730);
   U4448 : NBUFFX2 port map( INP => n4755, Z => n4729);
   U4449 : NBUFFX2 port map( INP => n4756, Z => n4725);
   U4450 : NBUFFX2 port map( INP => n4756, Z => n4727);
   U4451 : NBUFFX2 port map( INP => n4756, Z => n4726);
   U4452 : NBUFFX2 port map( INP => n4757, Z => n4722);
   U4453 : NBUFFX2 port map( INP => n4757, Z => n4724);
   U4454 : NBUFFX2 port map( INP => n4757, Z => n4723);
   U4455 : NBUFFX2 port map( INP => n4758, Z => n4719);
   U4456 : NBUFFX2 port map( INP => n4758, Z => n4721);
   U4457 : NBUFFX2 port map( INP => n4758, Z => n4720);
   U4458 : NBUFFX2 port map( INP => n4759, Z => n4716);
   U4459 : NBUFFX2 port map( INP => n4759, Z => n4718);
   U4460 : NBUFFX2 port map( INP => n4759, Z => n4717);
   U4461 : NBUFFX2 port map( INP => n4760, Z => n4713);
   U4462 : NBUFFX2 port map( INP => n4760, Z => n4715);
   U4463 : NBUFFX2 port map( INP => n4760, Z => n4714);
   U4464 : NBUFFX2 port map( INP => n4761, Z => n4710);
   U4465 : NBUFFX2 port map( INP => n4761, Z => n4712);
   U4466 : NBUFFX2 port map( INP => n4761, Z => n4711);
   U4467 : NBUFFX2 port map( INP => n4762, Z => n4707);
   U4468 : NBUFFX2 port map( INP => n4762, Z => n4709);
   U4469 : NBUFFX2 port map( INP => n4762, Z => n4708);
   U4470 : NBUFFX2 port map( INP => n4763, Z => n4704);
   U4471 : NBUFFX2 port map( INP => n4763, Z => n4706);
   U4472 : NBUFFX2 port map( INP => n4763, Z => n4705);
   U4473 : NBUFFX2 port map( INP => n4764, Z => n4701);
   U4474 : NBUFFX2 port map( INP => n4764, Z => n4703);
   U4475 : NBUFFX2 port map( INP => n4764, Z => n4702);
   U4476 : NBUFFX2 port map( INP => n4765, Z => n4698);
   U4477 : NBUFFX2 port map( INP => n4765, Z => n4700);
   U4478 : NBUFFX2 port map( INP => n4765, Z => n4699);
   U4479 : NBUFFX2 port map( INP => n4766, Z => n4695);
   U4480 : NBUFFX2 port map( INP => n4766, Z => n4697);
   U4481 : NBUFFX2 port map( INP => n4766, Z => n4696);
   U4482 : NBUFFX2 port map( INP => n4767, Z => n4692);
   U4483 : NBUFFX2 port map( INP => n4767, Z => n4693);
   U4484 : NBUFFX2 port map( INP => n4767, Z => n4694);
   U4485 : INVX0 port map( INP => RAMADDR2(2), ZN => n4514);
   U4486 : INVX0 port map( INP => RAMWRITE1, ZN => n5617);
   U4487 : NAND2X0 port map( IN1 => n33, IN2 => n23, QN => n32);
   U4488 : NAND2X0 port map( IN1 => n30, IN2 => n23, QN => n29);
   U4489 : NAND2X0 port map( IN1 => n22, IN2 => n23, QN => n21);
   U4490 : NBUFFX2 port map( INP => n4773, Z => n4750);
   U4491 : NBUFFX2 port map( INP => n4773, Z => n4751);
   U4492 : NBUFFX2 port map( INP => n4773, Z => n4752);
   U4493 : NBUFFX2 port map( INP => n4772, Z => n4753);
   U4494 : NBUFFX2 port map( INP => n4772, Z => n4754);
   U4495 : NBUFFX2 port map( INP => n4772, Z => n4755);
   U4496 : NBUFFX2 port map( INP => n4771, Z => n4756);
   U4497 : NBUFFX2 port map( INP => n4771, Z => n4757);
   U4498 : NBUFFX2 port map( INP => n4771, Z => n4758);
   U4499 : NBUFFX2 port map( INP => n4770, Z => n4759);
   U4500 : NBUFFX2 port map( INP => n4770, Z => n4760);
   U4501 : NBUFFX2 port map( INP => n4770, Z => n4761);
   U4502 : NBUFFX2 port map( INP => n4769, Z => n4762);
   U4503 : NBUFFX2 port map( INP => n4769, Z => n4763);
   U4504 : NBUFFX2 port map( INP => n4769, Z => n4764);
   U4505 : NBUFFX2 port map( INP => n4768, Z => n4765);
   U4506 : NBUFFX2 port map( INP => n4768, Z => n4766);
   U4507 : NBUFFX2 port map( INP => n4768, Z => n4767);
   U4508 : NBUFFX2 port map( INP => n4749, Z => n4746);
   U4509 : NBUFFX2 port map( INP => n4749, Z => n4748);
   U4510 : NBUFFX2 port map( INP => n4749, Z => n4747);
   U4511 : INVX0 port map( INP => RAMADDR2(0), ZN => n4515);
   U4512 : INVX0 port map( INP => RAMADDR2(3), ZN => n4513);
   U4513 : NOR2X0 port map( IN1 => n5616, IN2 => n2497, QN => n27);
   U4514 : NBUFFX2 port map( INP => clk, Z => n4773);
   U4515 : NBUFFX2 port map( INP => clk, Z => n4772);
   U4516 : NBUFFX2 port map( INP => clk, Z => n4771);
   U4517 : NBUFFX2 port map( INP => clk, Z => n4770);
   U4518 : NBUFFX2 port map( INP => clk, Z => n4769);
   U4519 : NBUFFX2 port map( INP => clk, Z => n4768);
   U4520 : NBUFFX2 port map( INP => n4774, Z => n4749);
   U4521 : NBUFFX2 port map( INP => clk, Z => n4774);
   U4522 : AOI221X1 port map( IN1 => RAM_0_3_port, IN2 => n2171, IN3 => 
                           RAM_1_3_port, IN4 => n3382, IN5 => n2841, QN => 
                           n3412);
   U4523 : AOI221X1 port map( IN1 => RAM_4_3_port, IN2 => n3407, IN3 => 
                           RAM_5_3_port, IN4 => n3401, IN5 => n2842, QN => 
                           n3411);
   U4524 : AO22X1 port map( IN1 => n5560, IN2 => RAMDIN1(66), IN3 => 
                           RAM_14_66_port, IN4 => n5542, Q => n241);
   U4525 : AO22X1 port map( IN1 => n5560, IN2 => RAMDIN1(67), IN3 => 
                           RAM_14_67_port, IN4 => n5542, Q => n242);
   U4526 : AOI221X1 port map( IN1 => RAM_4_102_port, IN2 => n3409, IN3 => 
                           RAM_5_102_port, IN4 => n3393, IN5 => n3238, QN => 
                           n3428);
   U4527 : AO22X1 port map( IN1 => n5558, IN2 => RAMDIN1(58), IN3 => 
                           RAM_14_58_port, IN4 => n5542, Q => n233);
   U4528 : AO22X1 port map( IN1 => n5560, IN2 => RAMDIN1(65), IN3 => 
                           RAM_14_65_port, IN4 => n5542, Q => n240);
   U4529 : AO22X1 port map( IN1 => n5559, IN2 => RAMDIN1(60), IN3 => 
                           RAM_14_60_port, IN4 => n5542, Q => n235);
   U4530 : AO22X1 port map( IN1 => n5560, IN2 => RAMDIN1(64), IN3 => 
                           RAM_14_64_port, IN4 => n5542, Q => n239);
   U4531 : AO22X1 port map( IN1 => n5558, IN2 => RAMDIN1(57), IN3 => 
                           RAM_14_57_port, IN4 => n5542, Q => n232);
   U4532 : AO22X1 port map( IN1 => n5559, IN2 => RAMDIN1(59), IN3 => 
                           RAM_14_59_port, IN4 => n5542, Q => n234);
   U4533 : AO22X1 port map( IN1 => n5559, IN2 => RAMDIN1(62), IN3 => 
                           RAM_14_62_port, IN4 => n5542, Q => n237);
   U4534 : AO22X1 port map( IN1 => n5559, IN2 => RAMDIN1(63), IN3 => 
                           RAM_14_63_port, IN4 => n5542, Q => n238);
   U4535 : AO22X1 port map( IN1 => n5558, IN2 => RAMDIN1(56), IN3 => 
                           RAM_14_56_port, IN4 => n5542, Q => n231);
   U4536 : AO22X1 port map( IN1 => n5559, IN2 => RAMDIN1(61), IN3 => 
                           RAM_14_61_port, IN4 => n5542, Q => n236);
   U4537 : AO22X1 port map( IN1 => RAMDIN1(58), IN2 => n5600, IN3 => 
                           RAM_15_58_port, IN4 => n5584, Q => n105);
   U4538 : AO22X1 port map( IN1 => n5600, IN2 => RAMDIN1(57), IN3 => 
                           RAM_15_57_port, IN4 => n5584, Q => n104);
   U4539 : AO22X1 port map( IN1 => RAMDIN1(56), IN2 => n5600, IN3 => 
                           RAM_15_56_port, IN4 => n5584, Q => n103);
   U4540 : NOR2X0 port map( IN1 => RAMADDR1(0), IN2 => RAMADDR1(1), QN => n2825
                           );
   U4541 : NOR2X0 port map( IN1 => n3359, IN2 => RAMADDR1(1), QN => n2826);
   U4542 : NOR2X0 port map( IN1 => RAMADDR1(2), IN2 => RAMADDR1(3), QN => n2823
                           );
   U4543 : NOR2X0 port map( IN1 => n3358, IN2 => RAMADDR1(3), QN => n2829);
   U4544 : AO22X1 port map( IN1 => RAM_7_0_port, IN2 => n2531, IN3 => 
                           RAM_6_0_port, IN4 => n2146, Q => n2830);
   U4545 : AO22X1 port map( IN1 => RAM_7_1_port, IN2 => n2514, IN3 => 
                           RAM_6_1_port, IN4 => n2148, Q => n2834);
   U4546 : AO22X1 port map( IN1 => RAM_7_2_port, IN2 => n2531, IN3 => 
                           RAM_6_2_port, IN4 => n2143, Q => n2838);
   U4547 : AO22X1 port map( IN1 => RAM_7_3_port, IN2 => n2530, IN3 => n2151, 
                           IN4 => RAM_6_3_port, Q => n2842);
   U4548 : AO22X1 port map( IN1 => RAM_15_4_port, IN2 => n3446, IN3 => 
                           RAM_14_4_port, IN4 => n2330, Q => n2844);
   U4549 : AO22X1 port map( IN1 => RAM_7_4_port, IN2 => n2517, IN3 => 
                           RAM_6_4_port, IN4 => n2149, Q => n2846);
   U4550 : AO22X1 port map( IN1 => RAM_15_5_port, IN2 => n3442, IN3 => 
                           RAM_14_5_port, IN4 => n2335, Q => n2848);
   U4551 : AO22X1 port map( IN1 => RAM_7_6_port, IN2 => n2521, IN3 => 
                           RAM_6_6_port, IN4 => n2140, Q => n2854);
   U4552 : AO22X1 port map( IN1 => RAM_7_7_port, IN2 => n2520, IN3 => 
                           RAM_6_7_port, IN4 => n2132, Q => n2858);
   U4553 : AO22X1 port map( IN1 => RAM_7_8_port, IN2 => n2522, IN3 => 
                           RAM_6_8_port, IN4 => n2134, Q => n2862);
   U4554 : AO22X1 port map( IN1 => RAM_7_12_port, IN2 => n2513, IN3 => 
                           RAM_6_12_port, IN4 => n2147, Q => n2878);
   U4555 : AO22X1 port map( IN1 => RAM_7_13_port, IN2 => n2528, IN3 => 
                           RAM_6_13_port, IN4 => n2139, Q => n2882);
   U4556 : AO22X1 port map( IN1 => RAM_7_14_port, IN2 => n2525, IN3 => 
                           RAM_6_14_port, IN4 => n2141, Q => n2886);
   U4557 : AO22X1 port map( IN1 => RAM_7_15_port, IN2 => n2524, IN3 => 
                           RAM_6_15_port, IN4 => n2149, Q => n2890);
   U4558 : AO22X1 port map( IN1 => RAM_7_16_port, IN2 => n2523, IN3 => 
                           RAM_6_16_port, IN4 => n2139, Q => n2894);
   U4559 : AO22X1 port map( IN1 => RAM_7_17_port, IN2 => n2522, IN3 => 
                           RAM_6_17_port, IN4 => n2143, Q => n2898);
   U4560 : AO22X1 port map( IN1 => RAM_7_18_port, IN2 => n2525, IN3 => 
                           RAM_6_18_port, IN4 => n2141, Q => n2902);
   U4561 : AO22X1 port map( IN1 => RAM_15_19_port, IN2 => n3446, IN3 => 
                           RAM_14_19_port, IN4 => n2322, Q => n2904);
   U4562 : AO22X1 port map( IN1 => RAM_7_21_port, IN2 => n2531, IN3 => 
                           RAM_6_21_port, IN4 => n2147, Q => n2914);
   U4563 : AO22X1 port map( IN1 => RAM_7_25_port, IN2 => n2513, IN3 => 
                           RAM_6_25_port, IN4 => n2144, Q => n2930);
   U4564 : AO22X1 port map( IN1 => RAM_7_26_port, IN2 => n2468, IN3 => 
                           RAM_6_26_port, IN4 => n2141, Q => n2934);
   U4565 : AO22X1 port map( IN1 => RAM_7_27_port, IN2 => n2530, IN3 => 
                           RAM_6_27_port, IN4 => n2140, Q => n2938);
   U4566 : AO22X1 port map( IN1 => RAM_7_28_port, IN2 => n2530, IN3 => 
                           RAM_6_28_port, IN4 => n2137, Q => n2942);
   U4567 : AO22X1 port map( IN1 => RAM_7_30_port, IN2 => n2518, IN3 => 
                           RAM_6_30_port, IN4 => n2133, Q => n2950);
   U4568 : AO22X1 port map( IN1 => RAM_7_31_port, IN2 => n2521, IN3 => 
                           RAM_6_31_port, IN4 => n2143, Q => n2954);
   U4569 : AO22X1 port map( IN1 => RAM_7_32_port, IN2 => n2518, IN3 => 
                           RAM_6_32_port, IN4 => n2149, Q => n2958);
   U4570 : AO22X1 port map( IN1 => RAM_7_34_port, IN2 => n2519, IN3 => 
                           RAM_6_34_port, IN4 => n2141, Q => n2966);
   U4571 : AO22X1 port map( IN1 => RAM_7_35_port, IN2 => n2527, IN3 => 
                           RAM_6_35_port, IN4 => n2143, Q => n2970);
   U4572 : AO22X1 port map( IN1 => RAM_7_37_port, IN2 => n2518, IN3 => 
                           RAM_6_37_port, IN4 => n2148, Q => n2978);
   U4573 : AO22X1 port map( IN1 => RAM_15_38_port, IN2 => n3436, IN3 => 
                           RAM_14_38_port, IN4 => n2321, Q => n2980);
   U4574 : AO22X1 port map( IN1 => RAM_7_40_port, IN2 => n2394, IN3 => 
                           RAM_6_40_port, IN4 => n2135, Q => n2990);
   U4575 : AO22X1 port map( IN1 => RAM_7_41_port, IN2 => n2340, IN3 => 
                           RAM_6_41_port, IN4 => n2152, Q => n2994);
   U4576 : AO22X1 port map( IN1 => RAM_7_42_port, IN2 => n2514, IN3 => 
                           RAM_6_42_port, IN4 => n2133, Q => n2998);
   U4577 : AO22X1 port map( IN1 => RAM_7_43_port, IN2 => n2340, IN3 => 
                           RAM_6_43_port, IN4 => n2138, Q => n3002);
   U4578 : AO22X1 port map( IN1 => RAM_7_44_port, IN2 => n2468, IN3 => 
                           RAM_6_44_port, IN4 => n2143, Q => n3006);
   U4579 : AO22X1 port map( IN1 => RAM_15_45_port, IN2 => n3439, IN3 => 
                           RAM_14_45_port, IN4 => n2339, Q => n3008);
   U4580 : AO22X1 port map( IN1 => RAM_7_46_port, IN2 => n2515, IN3 => 
                           RAM_6_46_port, IN4 => n2134, Q => n3014);
   U4581 : AO22X1 port map( IN1 => RAM_7_47_port, IN2 => n2517, IN3 => 
                           RAM_6_47_port, IN4 => n2134, Q => n3018);
   U4582 : AO22X1 port map( IN1 => RAM_7_48_port, IN2 => n2519, IN3 => 
                           RAM_6_48_port, IN4 => n2139, Q => n3022);
   U4583 : AO22X1 port map( IN1 => RAM_15_49_port, IN2 => n3442, IN3 => 
                           RAM_14_49_port, IN4 => n2337, Q => n3024);
   U4584 : AO22X1 port map( IN1 => RAM_7_49_port, IN2 => n2515, IN3 => 
                           RAM_6_49_port, IN4 => n2151, Q => n3026);
   U4585 : AO22X1 port map( IN1 => RAM_15_50_port, IN2 => n3433, IN3 => 
                           RAM_14_50_port, IN4 => n2336, Q => n3028);
   U4586 : AO22X1 port map( IN1 => RAM_7_50_port, IN2 => n2525, IN3 => 
                           RAM_6_50_port, IN4 => n2149, Q => n3030);
   U4587 : AO22X1 port map( IN1 => RAM_15_53_port, IN2 => n3446, IN3 => 
                           RAM_14_53_port, IN4 => n2320, Q => n3040);
   U4588 : AO22X1 port map( IN1 => RAM_7_53_port, IN2 => n2340, IN3 => 
                           RAM_6_53_port, IN4 => n2143, Q => n3042);
   U4589 : AO22X1 port map( IN1 => RAM_7_55_port, IN2 => n2530, IN3 => 
                           RAM_6_55_port, IN4 => n2151, Q => n3050);
   U4590 : AO22X1 port map( IN1 => RAM_15_56_port, IN2 => n3432, IN3 => 
                           RAM_14_56_port, IN4 => n2335, Q => n3052);
   U4591 : AO22X1 port map( IN1 => RAM_7_56_port, IN2 => n2531, IN3 => 
                           RAM_6_56_port, IN4 => n2142, Q => n3054);
   U4592 : AO22X1 port map( IN1 => RAM_7_58_port, IN2 => n2516, IN3 => 
                           RAM_6_58_port, IN4 => n2142, Q => n3062);
   U4593 : AO22X1 port map( IN1 => RAM_15_60_port, IN2 => n3437, IN3 => 
                           RAM_14_60_port, IN4 => n2323, Q => n3068);
   U4594 : AO22X1 port map( IN1 => RAM_7_61_port, IN2 => n2521, IN3 => 
                           RAM_6_61_port, IN4 => n2142, Q => n3074);
   U4595 : AO22X1 port map( IN1 => RAM_7_62_port, IN2 => n2513, IN3 => 
                           RAM_6_62_port, IN4 => n2132, Q => n3078);
   U4596 : AO22X1 port map( IN1 => RAM_15_65_port, IN2 => n3442, IN3 => 
                           RAM_14_65_port, IN4 => n2337, Q => n3088);
   U4597 : AO22X1 port map( IN1 => RAM_15_66_port, IN2 => n3444, IN3 => 
                           RAM_14_66_port, IN4 => n2337, Q => n3092);
   U4598 : AO22X1 port map( IN1 => RAM_7_66_port, IN2 => n2519, IN3 => 
                           RAM_6_66_port, IN4 => n2142, Q => n3094);
   U4599 : AO22X1 port map( IN1 => RAM_7_67_port, IN2 => n2523, IN3 => 
                           RAM_6_67_port, IN4 => n2145, Q => n3098);
   U4600 : AO22X1 port map( IN1 => RAM_15_68_port, IN2 => n3437, IN3 => 
                           RAM_14_68_port, IN4 => n2320, Q => n3100);
   U4601 : AO22X1 port map( IN1 => RAM_7_68_port, IN2 => n2517, IN3 => 
                           RAM_6_68_port, IN4 => n2134, Q => n3102);
   U4602 : AO22X1 port map( IN1 => RAM_7_69_port, IN2 => n2468, IN3 => 
                           RAM_6_69_port, IN4 => n2145, Q => n3106);
   U4603 : AO22X1 port map( IN1 => RAM_7_71_port, IN2 => n2528, IN3 => 
                           RAM_6_71_port, IN4 => n2144, Q => n3114);
   U4604 : AO22X1 port map( IN1 => RAM_7_72_port, IN2 => n2518, IN3 => 
                           RAM_6_72_port, IN4 => n2144, Q => n3118);
   U4605 : AO22X1 port map( IN1 => RAM_7_74_port, IN2 => n2340, IN3 => 
                           RAM_6_74_port, IN4 => n2146, Q => n3126);
   U4606 : AO22X1 port map( IN1 => RAM_7_76_port, IN2 => n2527, IN3 => 
                           RAM_6_76_port, IN4 => n2146, Q => n3134);
   U4607 : AO22X1 port map( IN1 => RAM_7_77_port, IN2 => n2529, IN3 => 
                           RAM_6_77_port, IN4 => n2146, Q => n3138);
   U4608 : AO22X1 port map( IN1 => RAM_7_78_port, IN2 => n2528, IN3 => 
                           RAM_6_78_port, IN4 => n2133, Q => n3142);
   U4609 : AO22X1 port map( IN1 => RAM_7_79_port, IN2 => n2528, IN3 => 
                           RAM_6_79_port, IN4 => n2137, Q => n3146);
   U4610 : AO22X1 port map( IN1 => RAM_7_80_port, IN2 => n2526, IN3 => 
                           RAM_6_80_port, IN4 => n2132, Q => n3150);
   U4611 : AO22X1 port map( IN1 => RAM_7_82_port, IN2 => n2517, IN3 => 
                           RAM_6_82_port, IN4 => n2138, Q => n3158);
   U4612 : AO22X1 port map( IN1 => RAM_7_84_port, IN2 => n2531, IN3 => 
                           RAM_6_84_port, IN4 => n2132, Q => n3166);
   U4613 : AO22X1 port map( IN1 => RAM_7_85_port, IN2 => n2525, IN3 => 
                           RAM_6_85_port, IN4 => n2150, Q => n3170);
   U4614 : AO22X1 port map( IN1 => RAM_15_86_port, IN2 => n3433, IN3 => 
                           RAM_14_86_port, IN4 => n2337, Q => n3172);
   U4615 : AO22X1 port map( IN1 => RAM_7_87_port, IN2 => n2529, IN3 => 
                           RAM_6_87_port, IN4 => n2136, Q => n3178);
   U4616 : AO22X1 port map( IN1 => RAM_7_88_port, IN2 => n2522, IN3 => 
                           RAM_6_88_port, IN4 => n2150, Q => n3182);
   U4617 : AO22X1 port map( IN1 => RAM_7_89_port, IN2 => n2529, IN3 => 
                           RAM_6_89_port, IN4 => n2144, Q => n3186);
   U4618 : AO22X1 port map( IN1 => RAM_7_91_port, IN2 => n2526, IN3 => 
                           RAM_6_91_port, IN4 => n2151, Q => n3194);
   U4619 : AO22X1 port map( IN1 => RAM_15_92_port, IN2 => n3434, IN3 => 
                           RAM_14_92_port, IN4 => n2322, Q => n3196);
   U4620 : AO22X1 port map( IN1 => RAM_7_92_port, IN2 => n2527, IN3 => 
                           RAM_6_92_port, IN4 => n2133, Q => n3198);
   U4621 : AO22X1 port map( IN1 => RAM_7_93_port, IN2 => n2524, IN3 => 
                           RAM_6_93_port, IN4 => n2134, Q => n3202);
   U4622 : AO22X1 port map( IN1 => RAM_15_94_port, IN2 => n3435, IN3 => 
                           RAM_14_94_port, IN4 => n2322, Q => n3204);
   U4623 : AO22X1 port map( IN1 => RAM_7_94_port, IN2 => n2513, IN3 => 
                           RAM_6_94_port, IN4 => n2132, Q => n3206);
   U4624 : AO22X1 port map( IN1 => RAM_7_96_port, IN2 => n2394, IN3 => 
                           RAM_6_96_port, IN4 => n2139, Q => n3214);
   U4625 : AO22X1 port map( IN1 => RAM_7_97_port, IN2 => n2520, IN3 => 
                           RAM_6_97_port, IN4 => n2148, Q => n3218);
   U4626 : AO22X1 port map( IN1 => RAM_7_100_port, IN2 => n2516, IN3 => n2142, 
                           IN4 => RAM_6_100_port, Q => n3230);
   U4627 : AO22X1 port map( IN1 => RAM_7_101_port, IN2 => n2523, IN3 => 
                           RAM_6_101_port, IN4 => n2136, Q => n3234);
   U4628 : AO22X1 port map( IN1 => RAM_7_103_port, IN2 => n2523, IN3 => 
                           RAM_6_103_port, IN4 => n2136, Q => n3242);
   U4629 : AO22X1 port map( IN1 => RAM_15_104_port, IN2 => n3432, IN3 => 
                           RAM_14_104_port, IN4 => n2326, Q => n3244);
   U4630 : AO22X1 port map( IN1 => RAM_7_104_port, IN2 => n2516, IN3 => 
                           RAM_6_104_port, IN4 => n2140, Q => n3246);
   U4631 : AO22X1 port map( IN1 => RAM_7_105_port, IN2 => n2518, IN3 => 
                           RAM_6_105_port, IN4 => n2145, Q => n3250);
   U4632 : AO22X1 port map( IN1 => RAM_7_106_port, IN2 => n2394, IN3 => 
                           RAM_6_106_port, IN4 => n2147, Q => n3254);
   U4633 : AO22X1 port map( IN1 => RAM_7_108_port, IN2 => n2468, IN3 => 
                           RAM_6_108_port, IN4 => n2150, Q => n3262);
   U4634 : AO22X1 port map( IN1 => RAM_7_109_port, IN2 => n2522, IN3 => 
                           RAM_6_109_port, IN4 => n2145, Q => n3266);
   U4635 : AO22X1 port map( IN1 => RAM_7_110_port, IN2 => n2515, IN3 => 
                           RAM_6_110_port, IN4 => n2145, Q => n3270);
   U4636 : AO221X1 port map( IN1 => RAM_8_112_port, IN2 => n3417, IN3 => 
                           RAM_9_112_port, IN4 => n3366, IN5 => n3275, Q => 
                           n3282);
   U4637 : AO221X1 port map( IN1 => RAM_0_112_port, IN2 => n2158, IN3 => 
                           RAM_1_112_port, IN4 => n3385, IN5 => n3277, Q => 
                           n3280);
   U4638 : AO22X1 port map( IN1 => RAM_7_112_port, IN2 => n2527, IN3 => 
                           RAM_6_112_port, IN4 => n2135, Q => n3278);
   U4639 : AO221X1 port map( IN1 => RAM_4_112_port, IN2 => n3404, IN3 => n3391,
                           IN4 => RAM_5_112_port, IN5 => n3278, Q => n3279);
   U4640 : AO22X1 port map( IN1 => RAM_7_114_port, IN2 => n2519, IN3 => 
                           RAM_6_114_port, IN4 => n2132, Q => n3290);
   U4641 : AO22X1 port map( IN1 => RAM_7_117_port, IN2 => n2520, IN3 => 
                           RAM_6_117_port, IN4 => n2146, Q => n3302);
   U4642 : AO22X1 port map( IN1 => RAM_15_118_port, IN2 => n3438, IN3 => 
                           RAM_14_118_port, IN4 => n2338, Q => n3304);
   U4643 : AO22X1 port map( IN1 => RAM_7_118_port, IN2 => n2514, IN3 => 
                           RAM_6_118_port, IN4 => n2146, Q => n3306);
   U4644 : AO22X1 port map( IN1 => RAM_7_119_port, IN2 => n2515, IN3 => 
                           RAM_6_119_port, IN4 => n2144, Q => n3310);
   U4645 : AO22X1 port map( IN1 => RAM_7_122_port, IN2 => n2526, IN3 => 
                           RAM_6_122_port, IN4 => n2174, Q => n3322);
   U4646 : AO22X1 port map( IN1 => RAM_7_123_port, IN2 => n2519, IN3 => 
                           RAM_6_123_port, IN4 => n2134, Q => n3326);
   U4647 : AO22X1 port map( IN1 => RAM_7_124_port, IN2 => n2529, IN3 => 
                           RAM_6_124_port, IN4 => n2135, Q => n3330);
   U4648 : AO22X1 port map( IN1 => RAM_7_126_port, IN2 => n2518, IN3 => 
                           RAM_6_126_port, IN4 => n2149, Q => n3338);
   U4649 : INVX0 port map( INP => RAMADDR1(0), ZN => n3359);
   U4650 : INVX0 port map( INP => RAMADDR1(2), ZN => n3358);
   U4651 : AOI221X1 port map( IN1 => RAM_12_3_port, IN2 => n2447, IN3 => 
                           RAM_13_3_port, IN4 => n3378, IN5 => n2840, QN => 
                           n3413);
   U4652 : NAND4X0 port map( IN1 => n3414, IN2 => n3413, IN3 => n3412, IN4 => 
                           n3411, QN => RAMDOUT1(3));
   U4653 : NBUFFX2 port map( INP => n3427, Z => n3415);
   U4654 : NBUFFX2 port map( INP => n3427, Z => n3416);
   U4655 : NBUFFX2 port map( INP => n3427, Z => n3417);
   U4656 : NBUFFX2 port map( INP => n3427, Z => n3418);
   U4657 : NBUFFX2 port map( INP => n3427, Z => n3419);
   U4658 : NBUFFX2 port map( INP => n3427, Z => n3420);
   U4659 : NBUFFX2 port map( INP => n3427, Z => n3423);
   U4660 : AOI221X1 port map( IN1 => RAM_8_102_port, IN2 => n3423, IN3 => 
                           RAM_9_102_port, IN4 => n2493, IN5 => n3235, QN => 
                           n3431);
   U4661 : NAND4X0 port map( IN1 => n3431, IN2 => n3430, IN3 => n3429, IN4 => 
                           n3428, QN => RAMDOUT1(102));
   U4662 : AOI221X1 port map( IN1 => RAM_0_102_port, IN2 => n2172, IN3 => 
                           RAM_1_102_port, IN4 => n3385, IN5 => n3237, QN => 
                           n3429);
   U4663 : AOI221X1 port map( IN1 => RAM_12_102_port, IN2 => n2451, IN3 => 
                           RAM_13_102_port, IN4 => n3379, IN5 => n3236, QN => 
                           n3430);
   U4664 : NBUFFX2 port map( INP => n3344, Z => n3439);
   U4665 : NBUFFX2 port map( INP => n3344, Z => n3440);
   U4666 : NBUFFX2 port map( INP => n3344, Z => n3441);
   U4667 : NBUFFX2 port map( INP => n3344, Z => n3446);
   U4668 : INVX0 port map( INP => n3464, ZN => n3449);
   U4669 : INVX0 port map( INP => n3464, ZN => n3450);
   U4670 : INVX0 port map( INP => n3464, ZN => n3452);
   U4671 : INVX0 port map( INP => n2499, ZN => n3455);
   U4672 : INVX0 port map( INP => n3463, ZN => n3456);
   U4673 : INVX0 port map( INP => n16, ZN => n3457);
   U4674 : INVX0 port map( INP => n3463, ZN => n3458);
   U4675 : INVX0 port map( INP => n2499, ZN => n3460);
   U4676 : INVX0 port map( INP => n3463, ZN => n3461);
   U4677 : INVX0 port map( INP => n3463, ZN => n3462);
   U4678 : INVX0 port map( INP => n3340, ZN => n3463);
   U4679 : NOR2X0 port map( IN1 => n4513, IN2 => RAMADDR2(2), QN => n3465);
   U4680 : NOR2X0 port map( IN1 => RAMADDR2(0), IN2 => RAMADDR2(1), QN => n3471
                           );
   U4681 : NOR2X0 port map( IN1 => n4515, IN2 => RAMADDR2(1), QN => n3472);
   U4682 : AND2X1 port map( IN1 => RAMADDR2(1), IN2 => RAMADDR2(0), Q => n3473)
                           ;
   U4683 : AND2X1 port map( IN1 => RAMADDR2(1), IN2 => n4515, Q => n3474);
   U4684 : AO22X1 port map( IN1 => RAM_11_0_port, IN2 => n4537, IN3 => 
                           RAM_10_0_port, IN4 => n4526, Q => n3466);
   U4685 : AO221X1 port map( IN1 => RAM_8_0_port, IN2 => n4559, IN3 => 
                           RAM_9_0_port, IN4 => n4548, IN5 => n3466, Q => n3480
                           );
   U4686 : NOR2X0 port map( IN1 => n4513, IN2 => n4514, QN => n3467);
   U4687 : AO22X1 port map( IN1 => RAM_15_0_port, IN2 => n4581, IN3 => 
                           RAM_14_0_port, IN4 => n4570, Q => n3468);
   U4688 : AO221X1 port map( IN1 => RAM_12_0_port, IN2 => n4603, IN3 => 
                           RAM_13_0_port, IN4 => n4592, IN5 => n3468, Q => 
                           n3479);
   U4689 : NOR2X0 port map( IN1 => RAMADDR2(2), IN2 => RAMADDR2(3), QN => n3469
                           );
   U4690 : AO22X1 port map( IN1 => RAM_3_0_port, IN2 => n4625, IN3 => 
                           RAM_2_0_port, IN4 => n4614, Q => n3470);
   U4691 : AO221X1 port map( IN1 => RAM_0_0_port, IN2 => n4647, IN3 => 
                           RAM_1_0_port, IN4 => n4636, IN5 => n3470, Q => n3478
                           );
   U4692 : NOR2X0 port map( IN1 => n4514, IN2 => RAMADDR2(3), QN => n3475);
   U4693 : AO22X1 port map( IN1 => RAM_7_0_port, IN2 => n4669, IN3 => 
                           RAM_6_0_port, IN4 => n4658, Q => n3476);
   U4694 : AO221X1 port map( IN1 => RAM_4_0_port, IN2 => n4691, IN3 => 
                           RAM_5_0_port, IN4 => n4680, IN5 => n3476, Q => n3477
                           );
   U4695 : OR4X1 port map( IN1 => n3480, IN2 => n3479, IN3 => n3478, IN4 => 
                           n3477, Q => RAMDOUT2(0));
   U4696 : AO22X1 port map( IN1 => RAM_11_1_port, IN2 => n4537, IN3 => 
                           RAM_10_1_port, IN4 => n4526, Q => n3481);
   U4697 : AO221X1 port map( IN1 => RAM_8_1_port, IN2 => n4559, IN3 => 
                           RAM_9_1_port, IN4 => n4548, IN5 => n3481, Q => n3488
                           );
   U4698 : AO22X1 port map( IN1 => RAM_15_1_port, IN2 => n4581, IN3 => 
                           RAM_14_1_port, IN4 => n4570, Q => n3482);
   U4699 : AO221X1 port map( IN1 => RAM_12_1_port, IN2 => n4603, IN3 => 
                           RAM_13_1_port, IN4 => n4592, IN5 => n3482, Q => 
                           n3487);
   U4700 : AO22X1 port map( IN1 => RAM_3_1_port, IN2 => n4625, IN3 => 
                           RAM_2_1_port, IN4 => n4614, Q => n3483);
   U4701 : AO221X1 port map( IN1 => RAM_0_1_port, IN2 => n4647, IN3 => 
                           RAM_1_1_port, IN4 => n4636, IN5 => n3483, Q => n3486
                           );
   U4702 : AO22X1 port map( IN1 => RAM_7_1_port, IN2 => n4669, IN3 => 
                           RAM_6_1_port, IN4 => n4658, Q => n3484);
   U4703 : AO221X1 port map( IN1 => RAM_4_1_port, IN2 => n4691, IN3 => 
                           RAM_5_1_port, IN4 => n4680, IN5 => n3484, Q => n3485
                           );
   U4704 : OR4X1 port map( IN1 => n3488, IN2 => n3487, IN3 => n3486, IN4 => 
                           n3485, Q => RAMDOUT2(1));
   U4705 : AO22X1 port map( IN1 => RAM_11_2_port, IN2 => n4537, IN3 => 
                           RAM_10_2_port, IN4 => n4526, Q => n3489);
   U4706 : AO221X1 port map( IN1 => RAM_8_2_port, IN2 => n4559, IN3 => 
                           RAM_9_2_port, IN4 => n4548, IN5 => n3489, Q => n3496
                           );
   U4707 : AO22X1 port map( IN1 => RAM_15_2_port, IN2 => n4581, IN3 => 
                           RAM_14_2_port, IN4 => n4570, Q => n3490);
   U4708 : AO221X1 port map( IN1 => RAM_12_2_port, IN2 => n4603, IN3 => 
                           RAM_13_2_port, IN4 => n4592, IN5 => n3490, Q => 
                           n3495);
   U4709 : AO22X1 port map( IN1 => RAM_3_2_port, IN2 => n4625, IN3 => 
                           RAM_2_2_port, IN4 => n4614, Q => n3491);
   U4710 : AO221X1 port map( IN1 => RAM_0_2_port, IN2 => n4647, IN3 => 
                           RAM_1_2_port, IN4 => n4636, IN5 => n3491, Q => n3494
                           );
   U4711 : AO22X1 port map( IN1 => RAM_7_2_port, IN2 => n4669, IN3 => 
                           RAM_6_2_port, IN4 => n4658, Q => n3492);
   U4712 : AO221X1 port map( IN1 => RAM_4_2_port, IN2 => n4691, IN3 => 
                           RAM_5_2_port, IN4 => n4680, IN5 => n3492, Q => n3493
                           );
   U4713 : OR4X1 port map( IN1 => n3496, IN2 => n3495, IN3 => n3494, IN4 => 
                           n3493, Q => RAMDOUT2(2));
   U4714 : AO22X1 port map( IN1 => RAM_11_3_port, IN2 => n4537, IN3 => 
                           RAM_10_3_port, IN4 => n4526, Q => n3497);
   U4715 : AO221X1 port map( IN1 => RAM_8_3_port, IN2 => n4559, IN3 => 
                           RAM_9_3_port, IN4 => n4548, IN5 => n3497, Q => n3504
                           );
   U4716 : AO22X1 port map( IN1 => RAM_15_3_port, IN2 => n4581, IN3 => 
                           RAM_14_3_port, IN4 => n4570, Q => n3498);
   U4717 : AO221X1 port map( IN1 => RAM_12_3_port, IN2 => n4603, IN3 => 
                           RAM_13_3_port, IN4 => n4592, IN5 => n3498, Q => 
                           n3503);
   U4718 : AO22X1 port map( IN1 => RAM_3_3_port, IN2 => n4625, IN3 => 
                           RAM_2_3_port, IN4 => n4614, Q => n3499);
   U4719 : AO221X1 port map( IN1 => RAM_0_3_port, IN2 => n4647, IN3 => 
                           RAM_1_3_port, IN4 => n4636, IN5 => n3499, Q => n3502
                           );
   U4720 : AO22X1 port map( IN1 => RAM_7_3_port, IN2 => n4669, IN3 => 
                           RAM_6_3_port, IN4 => n4658, Q => n3500);
   U4721 : AO221X1 port map( IN1 => RAM_4_3_port, IN2 => n4691, IN3 => 
                           RAM_5_3_port, IN4 => n4680, IN5 => n3500, Q => n3501
                           );
   U4722 : OR4X1 port map( IN1 => n3504, IN2 => n3503, IN3 => n3502, IN4 => 
                           n3501, Q => RAMDOUT2(3));
   U4723 : AO22X1 port map( IN1 => RAM_11_4_port, IN2 => n4537, IN3 => 
                           RAM_10_4_port, IN4 => n4526, Q => n3505);
   U4724 : AO221X1 port map( IN1 => RAM_8_4_port, IN2 => n4559, IN3 => 
                           RAM_9_4_port, IN4 => n4548, IN5 => n3505, Q => n3512
                           );
   U4725 : AO22X1 port map( IN1 => RAM_15_4_port, IN2 => n4581, IN3 => 
                           RAM_14_4_port, IN4 => n4570, Q => n3506);
   U4726 : AO221X1 port map( IN1 => RAM_12_4_port, IN2 => n4603, IN3 => 
                           RAM_13_4_port, IN4 => n4592, IN5 => n3506, Q => 
                           n3511);
   U4727 : AO22X1 port map( IN1 => RAM_3_4_port, IN2 => n4625, IN3 => 
                           RAM_2_4_port, IN4 => n4614, Q => n3507);
   U4728 : AO221X1 port map( IN1 => RAM_0_4_port, IN2 => n4647, IN3 => 
                           RAM_1_4_port, IN4 => n4636, IN5 => n3507, Q => n3510
                           );
   U4729 : AO22X1 port map( IN1 => RAM_7_4_port, IN2 => n4669, IN3 => 
                           RAM_6_4_port, IN4 => n4658, Q => n3508);
   U4730 : AO221X1 port map( IN1 => RAM_4_4_port, IN2 => n4691, IN3 => 
                           RAM_5_4_port, IN4 => n4680, IN5 => n3508, Q => n3509
                           );
   U4731 : OR4X1 port map( IN1 => n3512, IN2 => n3511, IN3 => n3510, IN4 => 
                           n3509, Q => RAMDOUT2(4));
   U4732 : AO22X1 port map( IN1 => RAM_11_5_port, IN2 => n4537, IN3 => 
                           RAM_10_5_port, IN4 => n4526, Q => n3513);
   U4733 : AO221X1 port map( IN1 => RAM_8_5_port, IN2 => n4559, IN3 => 
                           RAM_9_5_port, IN4 => n4548, IN5 => n3513, Q => n3520
                           );
   U4734 : AO22X1 port map( IN1 => RAM_15_5_port, IN2 => n4581, IN3 => 
                           RAM_14_5_port, IN4 => n4570, Q => n3514);
   U4735 : AO221X1 port map( IN1 => RAM_12_5_port, IN2 => n4603, IN3 => 
                           RAM_13_5_port, IN4 => n4592, IN5 => n3514, Q => 
                           n3519);
   U4736 : AO22X1 port map( IN1 => RAM_3_5_port, IN2 => n4625, IN3 => 
                           RAM_2_5_port, IN4 => n4614, Q => n3515);
   U4737 : AO221X1 port map( IN1 => RAM_0_5_port, IN2 => n4647, IN3 => 
                           RAM_1_5_port, IN4 => n4636, IN5 => n3515, Q => n3518
                           );
   U4738 : AO22X1 port map( IN1 => RAM_7_5_port, IN2 => n4669, IN3 => 
                           RAM_6_5_port, IN4 => n4658, Q => n3516);
   U4739 : AO221X1 port map( IN1 => RAM_4_5_port, IN2 => n4691, IN3 => 
                           RAM_5_5_port, IN4 => n4680, IN5 => n3516, Q => n3517
                           );
   U4740 : OR4X1 port map( IN1 => n3520, IN2 => n3519, IN3 => n3518, IN4 => 
                           n3517, Q => RAMDOUT2(5));
   U4741 : AO22X1 port map( IN1 => RAM_11_6_port, IN2 => n4537, IN3 => 
                           RAM_10_6_port, IN4 => n4526, Q => n3521);
   U4742 : AO221X1 port map( IN1 => RAM_8_6_port, IN2 => n4559, IN3 => 
                           RAM_9_6_port, IN4 => n4548, IN5 => n3521, Q => n3528
                           );
   U4743 : AO22X1 port map( IN1 => RAM_15_6_port, IN2 => n4581, IN3 => 
                           RAM_14_6_port, IN4 => n4570, Q => n3522);
   U4744 : AO221X1 port map( IN1 => RAM_12_6_port, IN2 => n4603, IN3 => 
                           RAM_13_6_port, IN4 => n4592, IN5 => n3522, Q => 
                           n3527);
   U4745 : AO22X1 port map( IN1 => RAM_3_6_port, IN2 => n4625, IN3 => 
                           RAM_2_6_port, IN4 => n4614, Q => n3523);
   U4746 : AO221X1 port map( IN1 => RAM_0_6_port, IN2 => n4647, IN3 => 
                           RAM_1_6_port, IN4 => n4636, IN5 => n3523, Q => n3526
                           );
   U4747 : AO22X1 port map( IN1 => RAM_7_6_port, IN2 => n4669, IN3 => 
                           RAM_6_6_port, IN4 => n4658, Q => n3524);
   U4748 : AO221X1 port map( IN1 => RAM_4_6_port, IN2 => n4691, IN3 => 
                           RAM_5_6_port, IN4 => n4680, IN5 => n3524, Q => n3525
                           );
   U4749 : OR4X1 port map( IN1 => n3528, IN2 => n3527, IN3 => n3526, IN4 => 
                           n3525, Q => RAMDOUT2(6));
   U4750 : AO22X1 port map( IN1 => RAM_11_7_port, IN2 => n4537, IN3 => 
                           RAM_10_7_port, IN4 => n4526, Q => n3529);
   U4751 : AO221X1 port map( IN1 => RAM_8_7_port, IN2 => n4559, IN3 => 
                           RAM_9_7_port, IN4 => n4548, IN5 => n3529, Q => n3536
                           );
   U4752 : AO22X1 port map( IN1 => RAM_15_7_port, IN2 => n4581, IN3 => 
                           RAM_14_7_port, IN4 => n4570, Q => n3530);
   U4753 : AO221X1 port map( IN1 => RAM_12_7_port, IN2 => n4603, IN3 => 
                           RAM_13_7_port, IN4 => n4592, IN5 => n3530, Q => 
                           n3535);
   U4754 : AO22X1 port map( IN1 => RAM_3_7_port, IN2 => n4625, IN3 => 
                           RAM_2_7_port, IN4 => n4614, Q => n3531);
   U4755 : AO221X1 port map( IN1 => RAM_0_7_port, IN2 => n4647, IN3 => 
                           RAM_1_7_port, IN4 => n4636, IN5 => n3531, Q => n3534
                           );
   U4756 : AO22X1 port map( IN1 => RAM_7_7_port, IN2 => n4669, IN3 => 
                           RAM_6_7_port, IN4 => n4658, Q => n3532);
   U4757 : AO221X1 port map( IN1 => RAM_4_7_port, IN2 => n4691, IN3 => 
                           RAM_5_7_port, IN4 => n4680, IN5 => n3532, Q => n3533
                           );
   U4758 : OR4X1 port map( IN1 => n3536, IN2 => n3535, IN3 => n3534, IN4 => 
                           n3533, Q => RAMDOUT2(7));
   U4759 : AO22X1 port map( IN1 => RAM_11_8_port, IN2 => n4537, IN3 => 
                           RAM_10_8_port, IN4 => n4526, Q => n3537);
   U4760 : AO221X1 port map( IN1 => RAM_8_8_port, IN2 => n4559, IN3 => 
                           RAM_9_8_port, IN4 => n4548, IN5 => n3537, Q => n3544
                           );
   U4761 : AO22X1 port map( IN1 => RAM_15_8_port, IN2 => n4581, IN3 => 
                           RAM_14_8_port, IN4 => n4570, Q => n3538);
   U4762 : AO221X1 port map( IN1 => RAM_12_8_port, IN2 => n4603, IN3 => 
                           RAM_13_8_port, IN4 => n4592, IN5 => n3538, Q => 
                           n3543);
   U4763 : AO22X1 port map( IN1 => RAM_3_8_port, IN2 => n4625, IN3 => 
                           RAM_2_8_port, IN4 => n4614, Q => n3539);
   U4764 : AO221X1 port map( IN1 => RAM_0_8_port, IN2 => n4647, IN3 => 
                           RAM_1_8_port, IN4 => n4636, IN5 => n3539, Q => n3542
                           );
   U4765 : AO22X1 port map( IN1 => RAM_7_8_port, IN2 => n4669, IN3 => 
                           RAM_6_8_port, IN4 => n4658, Q => n3540);
   U4766 : AO221X1 port map( IN1 => RAM_4_8_port, IN2 => n4691, IN3 => 
                           RAM_5_8_port, IN4 => n4680, IN5 => n3540, Q => n3541
                           );
   U4767 : OR4X1 port map( IN1 => n3544, IN2 => n3543, IN3 => n3542, IN4 => 
                           n3541, Q => RAMDOUT2(8));
   U4768 : AO22X1 port map( IN1 => RAM_11_9_port, IN2 => n4537, IN3 => 
                           RAM_10_9_port, IN4 => n4526, Q => n3545);
   U4769 : AO221X1 port map( IN1 => RAM_8_9_port, IN2 => n4559, IN3 => 
                           RAM_9_9_port, IN4 => n4548, IN5 => n3545, Q => n3552
                           );
   U4770 : AO22X1 port map( IN1 => RAM_15_9_port, IN2 => n4581, IN3 => 
                           RAM_14_9_port, IN4 => n4570, Q => n3546);
   U4771 : AO221X1 port map( IN1 => RAM_12_9_port, IN2 => n4603, IN3 => 
                           RAM_13_9_port, IN4 => n4592, IN5 => n3546, Q => 
                           n3551);
   U4772 : AO22X1 port map( IN1 => RAM_3_9_port, IN2 => n4625, IN3 => 
                           RAM_2_9_port, IN4 => n4614, Q => n3547);
   U4773 : AO221X1 port map( IN1 => RAM_0_9_port, IN2 => n4647, IN3 => 
                           RAM_1_9_port, IN4 => n4636, IN5 => n3547, Q => n3550
                           );
   U4774 : AO22X1 port map( IN1 => RAM_7_9_port, IN2 => n4669, IN3 => 
                           RAM_6_9_port, IN4 => n4658, Q => n3548);
   U4775 : AO221X1 port map( IN1 => RAM_4_9_port, IN2 => n4691, IN3 => 
                           RAM_5_9_port, IN4 => n4680, IN5 => n3548, Q => n3549
                           );
   U4776 : OR4X1 port map( IN1 => n3552, IN2 => n3551, IN3 => n3550, IN4 => 
                           n3549, Q => RAMDOUT2(9));
   U4777 : AO22X1 port map( IN1 => RAM_11_10_port, IN2 => n4537, IN3 => 
                           RAM_10_10_port, IN4 => n4526, Q => n3553);
   U4778 : AO221X1 port map( IN1 => RAM_8_10_port, IN2 => n4559, IN3 => 
                           RAM_9_10_port, IN4 => n4548, IN5 => n3553, Q => 
                           n3560);
   U4779 : AO22X1 port map( IN1 => RAM_15_10_port, IN2 => n4581, IN3 => 
                           RAM_14_10_port, IN4 => n4570, Q => n3554);
   U4780 : AO221X1 port map( IN1 => RAM_12_10_port, IN2 => n4603, IN3 => 
                           RAM_13_10_port, IN4 => n4592, IN5 => n3554, Q => 
                           n3559);
   U4781 : AO22X1 port map( IN1 => RAM_3_10_port, IN2 => n4625, IN3 => 
                           RAM_2_10_port, IN4 => n4614, Q => n3555);
   U4782 : AO221X1 port map( IN1 => RAM_0_10_port, IN2 => n4647, IN3 => 
                           RAM_1_10_port, IN4 => n4636, IN5 => n3555, Q => 
                           n3558);
   U4783 : AO22X1 port map( IN1 => RAM_7_10_port, IN2 => n4669, IN3 => 
                           RAM_6_10_port, IN4 => n4658, Q => n3556);
   U4784 : AO221X1 port map( IN1 => RAM_4_10_port, IN2 => n4691, IN3 => 
                           RAM_5_10_port, IN4 => n4680, IN5 => n3556, Q => 
                           n3557);
   U4785 : OR4X1 port map( IN1 => n3560, IN2 => n3559, IN3 => n3558, IN4 => 
                           n3557, Q => RAMDOUT2(10));
   U4786 : AO22X1 port map( IN1 => RAM_11_11_port, IN2 => n4537, IN3 => 
                           RAM_10_11_port, IN4 => n4526, Q => n3561);
   U4787 : AO221X1 port map( IN1 => RAM_8_11_port, IN2 => n4559, IN3 => 
                           RAM_9_11_port, IN4 => n4548, IN5 => n3561, Q => 
                           n3568);
   U4788 : AO22X1 port map( IN1 => RAM_15_11_port, IN2 => n4581, IN3 => 
                           RAM_14_11_port, IN4 => n4570, Q => n3562);
   U4789 : AO221X1 port map( IN1 => RAM_12_11_port, IN2 => n4603, IN3 => 
                           RAM_13_11_port, IN4 => n4592, IN5 => n3562, Q => 
                           n3567);
   U4790 : AO22X1 port map( IN1 => RAM_3_11_port, IN2 => n4625, IN3 => 
                           RAM_2_11_port, IN4 => n4614, Q => n3563);
   U4791 : AO221X1 port map( IN1 => RAM_0_11_port, IN2 => n4647, IN3 => 
                           RAM_1_11_port, IN4 => n4636, IN5 => n3563, Q => 
                           n3566);
   U4792 : AO22X1 port map( IN1 => RAM_7_11_port, IN2 => n4669, IN3 => 
                           RAM_6_11_port, IN4 => n4658, Q => n3564);
   U4793 : AO221X1 port map( IN1 => RAM_4_11_port, IN2 => n4691, IN3 => 
                           RAM_5_11_port, IN4 => n4680, IN5 => n3564, Q => 
                           n3565);
   U4794 : OR4X1 port map( IN1 => n3568, IN2 => n3567, IN3 => n3566, IN4 => 
                           n3565, Q => RAMDOUT2(11));
   U4795 : AO22X1 port map( IN1 => RAM_11_12_port, IN2 => n4536, IN3 => 
                           RAM_10_12_port, IN4 => n4525, Q => n3569);
   U4796 : AO221X1 port map( IN1 => RAM_8_12_port, IN2 => n4558, IN3 => 
                           RAM_9_12_port, IN4 => n4547, IN5 => n3569, Q => 
                           n3576);
   U4797 : AO22X1 port map( IN1 => RAM_15_12_port, IN2 => n4580, IN3 => 
                           RAM_14_12_port, IN4 => n4569, Q => n3570);
   U4798 : AO221X1 port map( IN1 => RAM_12_12_port, IN2 => n4602, IN3 => 
                           RAM_13_12_port, IN4 => n4591, IN5 => n3570, Q => 
                           n3575);
   U4799 : AO22X1 port map( IN1 => RAM_3_12_port, IN2 => n4624, IN3 => 
                           RAM_2_12_port, IN4 => n4613, Q => n3571);
   U4800 : AO221X1 port map( IN1 => RAM_0_12_port, IN2 => n4646, IN3 => 
                           RAM_1_12_port, IN4 => n4635, IN5 => n3571, Q => 
                           n3574);
   U4801 : AO22X1 port map( IN1 => RAM_7_12_port, IN2 => n4668, IN3 => 
                           RAM_6_12_port, IN4 => n4657, Q => n3572);
   U4802 : AO221X1 port map( IN1 => RAM_4_12_port, IN2 => n4690, IN3 => 
                           RAM_5_12_port, IN4 => n4679, IN5 => n3572, Q => 
                           n3573);
   U4803 : OR4X1 port map( IN1 => n3576, IN2 => n3575, IN3 => n3574, IN4 => 
                           n3573, Q => RAMDOUT2(12));
   U4804 : AO22X1 port map( IN1 => RAM_11_13_port, IN2 => n4536, IN3 => 
                           RAM_10_13_port, IN4 => n4525, Q => n3577);
   U4805 : AO221X1 port map( IN1 => RAM_8_13_port, IN2 => n4558, IN3 => 
                           RAM_9_13_port, IN4 => n4547, IN5 => n3577, Q => 
                           n3584);
   U4806 : AO22X1 port map( IN1 => RAM_15_13_port, IN2 => n4580, IN3 => 
                           RAM_14_13_port, IN4 => n4569, Q => n3578);
   U4807 : AO221X1 port map( IN1 => RAM_12_13_port, IN2 => n4602, IN3 => 
                           RAM_13_13_port, IN4 => n4591, IN5 => n3578, Q => 
                           n3583);
   U4808 : AO22X1 port map( IN1 => RAM_3_13_port, IN2 => n4624, IN3 => 
                           RAM_2_13_port, IN4 => n4613, Q => n3579);
   U4809 : AO221X1 port map( IN1 => RAM_0_13_port, IN2 => n4646, IN3 => 
                           RAM_1_13_port, IN4 => n4635, IN5 => n3579, Q => 
                           n3582);
   U4810 : AO22X1 port map( IN1 => RAM_7_13_port, IN2 => n4668, IN3 => 
                           RAM_6_13_port, IN4 => n4657, Q => n3580);
   U4811 : AO221X1 port map( IN1 => RAM_4_13_port, IN2 => n4690, IN3 => 
                           RAM_5_13_port, IN4 => n4679, IN5 => n3580, Q => 
                           n3581);
   U4812 : OR4X1 port map( IN1 => n3584, IN2 => n3583, IN3 => n3582, IN4 => 
                           n3581, Q => RAMDOUT2(13));
   U4813 : AO22X1 port map( IN1 => RAM_11_14_port, IN2 => n4536, IN3 => 
                           RAM_10_14_port, IN4 => n4525, Q => n3585);
   U4814 : AO221X1 port map( IN1 => RAM_8_14_port, IN2 => n4558, IN3 => 
                           RAM_9_14_port, IN4 => n4547, IN5 => n3585, Q => 
                           n3592);
   U4815 : AO22X1 port map( IN1 => RAM_15_14_port, IN2 => n4580, IN3 => 
                           RAM_14_14_port, IN4 => n4569, Q => n3586);
   U4816 : AO221X1 port map( IN1 => RAM_12_14_port, IN2 => n4602, IN3 => 
                           RAM_13_14_port, IN4 => n4591, IN5 => n3586, Q => 
                           n3591);
   U4817 : AO22X1 port map( IN1 => RAM_3_14_port, IN2 => n4624, IN3 => 
                           RAM_2_14_port, IN4 => n4613, Q => n3587);
   U4818 : AO221X1 port map( IN1 => RAM_0_14_port, IN2 => n4646, IN3 => 
                           RAM_1_14_port, IN4 => n4635, IN5 => n3587, Q => 
                           n3590);
   U4819 : AO22X1 port map( IN1 => RAM_7_14_port, IN2 => n4668, IN3 => 
                           RAM_6_14_port, IN4 => n4657, Q => n3588);
   U4820 : AO221X1 port map( IN1 => RAM_4_14_port, IN2 => n4690, IN3 => 
                           RAM_5_14_port, IN4 => n4679, IN5 => n3588, Q => 
                           n3589);
   U4821 : OR4X1 port map( IN1 => n3592, IN2 => n3591, IN3 => n3590, IN4 => 
                           n3589, Q => RAMDOUT2(14));
   U4822 : AO22X1 port map( IN1 => RAM_11_15_port, IN2 => n4536, IN3 => 
                           RAM_10_15_port, IN4 => n4525, Q => n3593);
   U4823 : AO221X1 port map( IN1 => RAM_8_15_port, IN2 => n4558, IN3 => 
                           RAM_9_15_port, IN4 => n4547, IN5 => n3593, Q => 
                           n3600);
   U4824 : AO22X1 port map( IN1 => RAM_15_15_port, IN2 => n4580, IN3 => 
                           RAM_14_15_port, IN4 => n4569, Q => n3594);
   U4825 : AO221X1 port map( IN1 => RAM_12_15_port, IN2 => n4602, IN3 => 
                           RAM_13_15_port, IN4 => n4591, IN5 => n3594, Q => 
                           n3599);
   U4826 : AO22X1 port map( IN1 => RAM_3_15_port, IN2 => n4624, IN3 => 
                           RAM_2_15_port, IN4 => n4613, Q => n3595);
   U4827 : AO221X1 port map( IN1 => RAM_0_15_port, IN2 => n4646, IN3 => 
                           RAM_1_15_port, IN4 => n4635, IN5 => n3595, Q => 
                           n3598);
   U4828 : AO22X1 port map( IN1 => RAM_7_15_port, IN2 => n4668, IN3 => 
                           RAM_6_15_port, IN4 => n4657, Q => n3596);
   U4829 : AO221X1 port map( IN1 => RAM_4_15_port, IN2 => n4690, IN3 => 
                           RAM_5_15_port, IN4 => n4679, IN5 => n3596, Q => 
                           n3597);
   U4830 : OR4X1 port map( IN1 => n3600, IN2 => n3599, IN3 => n3598, IN4 => 
                           n3597, Q => RAMDOUT2(15));
   U4831 : AO22X1 port map( IN1 => RAM_11_16_port, IN2 => n4536, IN3 => 
                           RAM_10_16_port, IN4 => n4525, Q => n3601);
   U4832 : AO221X1 port map( IN1 => RAM_8_16_port, IN2 => n4558, IN3 => 
                           RAM_9_16_port, IN4 => n4547, IN5 => n3601, Q => 
                           n3608);
   U4833 : AO22X1 port map( IN1 => RAM_15_16_port, IN2 => n4580, IN3 => 
                           RAM_14_16_port, IN4 => n4569, Q => n3602);
   U4834 : AO221X1 port map( IN1 => RAM_12_16_port, IN2 => n4602, IN3 => 
                           RAM_13_16_port, IN4 => n4591, IN5 => n3602, Q => 
                           n3607);
   U4835 : AO22X1 port map( IN1 => RAM_3_16_port, IN2 => n4624, IN3 => 
                           RAM_2_16_port, IN4 => n4613, Q => n3603);
   U4836 : AO221X1 port map( IN1 => RAM_0_16_port, IN2 => n4646, IN3 => 
                           RAM_1_16_port, IN4 => n4635, IN5 => n3603, Q => 
                           n3606);
   U4837 : AO22X1 port map( IN1 => RAM_7_16_port, IN2 => n4668, IN3 => 
                           RAM_6_16_port, IN4 => n4657, Q => n3604);
   U4838 : AO221X1 port map( IN1 => RAM_4_16_port, IN2 => n4690, IN3 => 
                           RAM_5_16_port, IN4 => n4679, IN5 => n3604, Q => 
                           n3605);
   U4839 : OR4X1 port map( IN1 => n3608, IN2 => n3607, IN3 => n3606, IN4 => 
                           n3605, Q => RAMDOUT2(16));
   U4840 : AO22X1 port map( IN1 => RAM_11_17_port, IN2 => n4536, IN3 => 
                           RAM_10_17_port, IN4 => n4525, Q => n3609);
   U4841 : AO221X1 port map( IN1 => RAM_8_17_port, IN2 => n4558, IN3 => 
                           RAM_9_17_port, IN4 => n4547, IN5 => n3609, Q => 
                           n3616);
   U4842 : AO22X1 port map( IN1 => RAM_15_17_port, IN2 => n4580, IN3 => 
                           RAM_14_17_port, IN4 => n4569, Q => n3610);
   U4843 : AO221X1 port map( IN1 => RAM_12_17_port, IN2 => n4602, IN3 => 
                           RAM_13_17_port, IN4 => n4591, IN5 => n3610, Q => 
                           n3615);
   U4844 : AO22X1 port map( IN1 => RAM_3_17_port, IN2 => n4624, IN3 => 
                           RAM_2_17_port, IN4 => n4613, Q => n3611);
   U4845 : AO221X1 port map( IN1 => RAM_0_17_port, IN2 => n4646, IN3 => 
                           RAM_1_17_port, IN4 => n4635, IN5 => n3611, Q => 
                           n3614);
   U4846 : AO22X1 port map( IN1 => RAM_7_17_port, IN2 => n4668, IN3 => 
                           RAM_6_17_port, IN4 => n4657, Q => n3612);
   U4847 : AO221X1 port map( IN1 => RAM_4_17_port, IN2 => n4690, IN3 => 
                           RAM_5_17_port, IN4 => n4679, IN5 => n3612, Q => 
                           n3613);
   U4848 : OR4X1 port map( IN1 => n3616, IN2 => n3615, IN3 => n3614, IN4 => 
                           n3613, Q => RAMDOUT2(17));
   U4849 : AO22X1 port map( IN1 => RAM_11_18_port, IN2 => n4536, IN3 => 
                           RAM_10_18_port, IN4 => n4525, Q => n3617);
   U4850 : AO221X1 port map( IN1 => RAM_8_18_port, IN2 => n4558, IN3 => 
                           RAM_9_18_port, IN4 => n4547, IN5 => n3617, Q => 
                           n3624);
   U4851 : AO22X1 port map( IN1 => RAM_15_18_port, IN2 => n4580, IN3 => 
                           RAM_14_18_port, IN4 => n4569, Q => n3618);
   U4852 : AO221X1 port map( IN1 => RAM_12_18_port, IN2 => n4602, IN3 => 
                           RAM_13_18_port, IN4 => n4591, IN5 => n3618, Q => 
                           n3623);
   U4853 : AO22X1 port map( IN1 => RAM_3_18_port, IN2 => n4624, IN3 => 
                           RAM_2_18_port, IN4 => n4613, Q => n3619);
   U4854 : AO221X1 port map( IN1 => RAM_0_18_port, IN2 => n4646, IN3 => 
                           RAM_1_18_port, IN4 => n4635, IN5 => n3619, Q => 
                           n3622);
   U4855 : AO22X1 port map( IN1 => RAM_7_18_port, IN2 => n4668, IN3 => 
                           RAM_6_18_port, IN4 => n4657, Q => n3620);
   U4856 : AO221X1 port map( IN1 => RAM_4_18_port, IN2 => n4690, IN3 => 
                           RAM_5_18_port, IN4 => n4679, IN5 => n3620, Q => 
                           n3621);
   U4857 : OR4X1 port map( IN1 => n3624, IN2 => n3623, IN3 => n3622, IN4 => 
                           n3621, Q => RAMDOUT2(18));
   U4858 : AO22X1 port map( IN1 => RAM_11_19_port, IN2 => n4536, IN3 => 
                           RAM_10_19_port, IN4 => n4525, Q => n3625);
   U4859 : AO221X1 port map( IN1 => RAM_8_19_port, IN2 => n4558, IN3 => 
                           RAM_9_19_port, IN4 => n4547, IN5 => n3625, Q => 
                           n3632);
   U4860 : AO22X1 port map( IN1 => RAM_15_19_port, IN2 => n4580, IN3 => 
                           RAM_14_19_port, IN4 => n4569, Q => n3626);
   U4861 : AO221X1 port map( IN1 => RAM_12_19_port, IN2 => n4602, IN3 => 
                           RAM_13_19_port, IN4 => n4591, IN5 => n3626, Q => 
                           n3631);
   U4862 : AO22X1 port map( IN1 => RAM_3_19_port, IN2 => n4624, IN3 => 
                           RAM_2_19_port, IN4 => n4613, Q => n3627);
   U4863 : AO221X1 port map( IN1 => RAM_0_19_port, IN2 => n4646, IN3 => 
                           RAM_1_19_port, IN4 => n4635, IN5 => n3627, Q => 
                           n3630);
   U4864 : AO22X1 port map( IN1 => RAM_7_19_port, IN2 => n4668, IN3 => 
                           RAM_6_19_port, IN4 => n4657, Q => n3628);
   U4865 : AO221X1 port map( IN1 => RAM_4_19_port, IN2 => n4690, IN3 => 
                           RAM_5_19_port, IN4 => n4679, IN5 => n3628, Q => 
                           n3629);
   U4866 : OR4X1 port map( IN1 => n3632, IN2 => n3631, IN3 => n3630, IN4 => 
                           n3629, Q => RAMDOUT2(19));
   U4867 : AO22X1 port map( IN1 => RAM_11_20_port, IN2 => n4536, IN3 => 
                           RAM_10_20_port, IN4 => n4525, Q => n3633);
   U4868 : AO221X1 port map( IN1 => RAM_8_20_port, IN2 => n4558, IN3 => 
                           RAM_9_20_port, IN4 => n4547, IN5 => n3633, Q => 
                           n3640);
   U4869 : AO22X1 port map( IN1 => RAM_15_20_port, IN2 => n4580, IN3 => 
                           RAM_14_20_port, IN4 => n4569, Q => n3634);
   U4870 : AO221X1 port map( IN1 => RAM_12_20_port, IN2 => n4602, IN3 => 
                           RAM_13_20_port, IN4 => n4591, IN5 => n3634, Q => 
                           n3639);
   U4871 : AO22X1 port map( IN1 => RAM_3_20_port, IN2 => n4624, IN3 => 
                           RAM_2_20_port, IN4 => n4613, Q => n3635);
   U4872 : AO221X1 port map( IN1 => RAM_0_20_port, IN2 => n4646, IN3 => 
                           RAM_1_20_port, IN4 => n4635, IN5 => n3635, Q => 
                           n3638);
   U4873 : AO22X1 port map( IN1 => RAM_7_20_port, IN2 => n4668, IN3 => 
                           RAM_6_20_port, IN4 => n4657, Q => n3636);
   U4874 : AO221X1 port map( IN1 => RAM_4_20_port, IN2 => n4690, IN3 => 
                           RAM_5_20_port, IN4 => n4679, IN5 => n3636, Q => 
                           n3637);
   U4875 : OR4X1 port map( IN1 => n3640, IN2 => n3639, IN3 => n3638, IN4 => 
                           n3637, Q => RAMDOUT2(20));
   U4876 : AO22X1 port map( IN1 => RAM_11_21_port, IN2 => n4536, IN3 => 
                           RAM_10_21_port, IN4 => n4525, Q => n3641);
   U4877 : AO221X1 port map( IN1 => RAM_8_21_port, IN2 => n4558, IN3 => 
                           RAM_9_21_port, IN4 => n4547, IN5 => n3641, Q => 
                           n3648);
   U4878 : AO22X1 port map( IN1 => RAM_15_21_port, IN2 => n4580, IN3 => 
                           RAM_14_21_port, IN4 => n4569, Q => n3642);
   U4879 : AO221X1 port map( IN1 => RAM_12_21_port, IN2 => n4602, IN3 => 
                           RAM_13_21_port, IN4 => n4591, IN5 => n3642, Q => 
                           n3647);
   U4880 : AO22X1 port map( IN1 => RAM_3_21_port, IN2 => n4624, IN3 => 
                           RAM_2_21_port, IN4 => n4613, Q => n3643);
   U4881 : AO221X1 port map( IN1 => RAM_0_21_port, IN2 => n4646, IN3 => 
                           RAM_1_21_port, IN4 => n4635, IN5 => n3643, Q => 
                           n3646);
   U4882 : AO22X1 port map( IN1 => RAM_7_21_port, IN2 => n4668, IN3 => 
                           RAM_6_21_port, IN4 => n4657, Q => n3644);
   U4883 : AO221X1 port map( IN1 => RAM_4_21_port, IN2 => n4690, IN3 => 
                           RAM_5_21_port, IN4 => n4679, IN5 => n3644, Q => 
                           n3645);
   U4884 : OR4X1 port map( IN1 => n3648, IN2 => n3647, IN3 => n3646, IN4 => 
                           n3645, Q => RAMDOUT2(21));
   U4885 : AO22X1 port map( IN1 => RAM_11_22_port, IN2 => n4536, IN3 => 
                           RAM_10_22_port, IN4 => n4525, Q => n3649);
   U4886 : AO221X1 port map( IN1 => RAM_8_22_port, IN2 => n4558, IN3 => 
                           RAM_9_22_port, IN4 => n4547, IN5 => n3649, Q => 
                           n3656);
   U4887 : AO22X1 port map( IN1 => RAM_15_22_port, IN2 => n4580, IN3 => 
                           RAM_14_22_port, IN4 => n4569, Q => n3650);
   U4888 : AO221X1 port map( IN1 => RAM_12_22_port, IN2 => n4602, IN3 => 
                           RAM_13_22_port, IN4 => n4591, IN5 => n3650, Q => 
                           n3655);
   U4889 : AO22X1 port map( IN1 => RAM_3_22_port, IN2 => n4624, IN3 => 
                           RAM_2_22_port, IN4 => n4613, Q => n3651);
   U4890 : AO221X1 port map( IN1 => RAM_0_22_port, IN2 => n4646, IN3 => 
                           RAM_1_22_port, IN4 => n4635, IN5 => n3651, Q => 
                           n3654);
   U4891 : AO22X1 port map( IN1 => RAM_7_22_port, IN2 => n4668, IN3 => 
                           RAM_6_22_port, IN4 => n4657, Q => n3652);
   U4892 : AO221X1 port map( IN1 => RAM_4_22_port, IN2 => n4690, IN3 => 
                           RAM_5_22_port, IN4 => n4679, IN5 => n3652, Q => 
                           n3653);
   U4893 : OR4X1 port map( IN1 => n3656, IN2 => n3655, IN3 => n3654, IN4 => 
                           n3653, Q => RAMDOUT2(22));
   U4894 : AO22X1 port map( IN1 => RAM_11_23_port, IN2 => n4536, IN3 => 
                           RAM_10_23_port, IN4 => n4525, Q => n3657);
   U4895 : AO221X1 port map( IN1 => RAM_8_23_port, IN2 => n4558, IN3 => 
                           RAM_9_23_port, IN4 => n4547, IN5 => n3657, Q => 
                           n3664);
   U4896 : AO22X1 port map( IN1 => RAM_15_23_port, IN2 => n4580, IN3 => 
                           RAM_14_23_port, IN4 => n4569, Q => n3658);
   U4897 : AO221X1 port map( IN1 => RAM_12_23_port, IN2 => n4602, IN3 => 
                           RAM_13_23_port, IN4 => n4591, IN5 => n3658, Q => 
                           n3663);
   U4898 : AO22X1 port map( IN1 => RAM_3_23_port, IN2 => n4624, IN3 => 
                           RAM_2_23_port, IN4 => n4613, Q => n3659);
   U4899 : AO221X1 port map( IN1 => RAM_0_23_port, IN2 => n4646, IN3 => 
                           RAM_1_23_port, IN4 => n4635, IN5 => n3659, Q => 
                           n3662);
   U4900 : AO22X1 port map( IN1 => RAM_7_23_port, IN2 => n4668, IN3 => 
                           RAM_6_23_port, IN4 => n4657, Q => n3660);
   U4901 : AO221X1 port map( IN1 => RAM_4_23_port, IN2 => n4690, IN3 => 
                           RAM_5_23_port, IN4 => n4679, IN5 => n3660, Q => 
                           n3661);
   U4902 : OR4X1 port map( IN1 => n3664, IN2 => n3663, IN3 => n3662, IN4 => 
                           n3661, Q => RAMDOUT2(23));
   U4903 : AO22X1 port map( IN1 => RAM_11_24_port, IN2 => n4535, IN3 => 
                           RAM_10_24_port, IN4 => n4524, Q => n3665);
   U4904 : AO221X1 port map( IN1 => RAM_8_24_port, IN2 => n4557, IN3 => 
                           RAM_9_24_port, IN4 => n4546, IN5 => n3665, Q => 
                           n3672);
   U4905 : AO22X1 port map( IN1 => RAM_15_24_port, IN2 => n4579, IN3 => 
                           RAM_14_24_port, IN4 => n4568, Q => n3666);
   U4906 : AO221X1 port map( IN1 => RAM_12_24_port, IN2 => n4601, IN3 => 
                           RAM_13_24_port, IN4 => n4590, IN5 => n3666, Q => 
                           n3671);
   U4907 : AO22X1 port map( IN1 => RAM_3_24_port, IN2 => n4623, IN3 => 
                           RAM_2_24_port, IN4 => n4612, Q => n3667);
   U4908 : AO221X1 port map( IN1 => RAM_0_24_port, IN2 => n4645, IN3 => 
                           RAM_1_24_port, IN4 => n4634, IN5 => n3667, Q => 
                           n3670);
   U4909 : AO22X1 port map( IN1 => RAM_7_24_port, IN2 => n4667, IN3 => 
                           RAM_6_24_port, IN4 => n4656, Q => n3668);
   U4910 : AO221X1 port map( IN1 => RAM_4_24_port, IN2 => n4689, IN3 => 
                           RAM_5_24_port, IN4 => n4678, IN5 => n3668, Q => 
                           n3669);
   U4911 : OR4X1 port map( IN1 => n3672, IN2 => n3671, IN3 => n3670, IN4 => 
                           n3669, Q => RAMDOUT2(24));
   U4912 : AO22X1 port map( IN1 => RAM_11_25_port, IN2 => n4535, IN3 => 
                           RAM_10_25_port, IN4 => n4524, Q => n3673);
   U4913 : AO221X1 port map( IN1 => RAM_8_25_port, IN2 => n4557, IN3 => 
                           RAM_9_25_port, IN4 => n4546, IN5 => n3673, Q => 
                           n3680);
   U4914 : AO22X1 port map( IN1 => RAM_15_25_port, IN2 => n4579, IN3 => 
                           RAM_14_25_port, IN4 => n4568, Q => n3674);
   U4915 : AO221X1 port map( IN1 => RAM_12_25_port, IN2 => n4601, IN3 => 
                           RAM_13_25_port, IN4 => n4590, IN5 => n3674, Q => 
                           n3679);
   U4916 : AO22X1 port map( IN1 => RAM_3_25_port, IN2 => n4623, IN3 => 
                           RAM_2_25_port, IN4 => n4612, Q => n3675);
   U4917 : AO221X1 port map( IN1 => RAM_0_25_port, IN2 => n4645, IN3 => 
                           RAM_1_25_port, IN4 => n4634, IN5 => n3675, Q => 
                           n3678);
   U4918 : AO22X1 port map( IN1 => RAM_7_25_port, IN2 => n4667, IN3 => 
                           RAM_6_25_port, IN4 => n4656, Q => n3676);
   U4919 : AO221X1 port map( IN1 => RAM_4_25_port, IN2 => n4689, IN3 => 
                           RAM_5_25_port, IN4 => n4678, IN5 => n3676, Q => 
                           n3677);
   U4920 : OR4X1 port map( IN1 => n3680, IN2 => n3679, IN3 => n3678, IN4 => 
                           n3677, Q => RAMDOUT2(25));
   U4921 : AO22X1 port map( IN1 => RAM_11_26_port, IN2 => n4535, IN3 => 
                           RAM_10_26_port, IN4 => n4524, Q => n3681);
   U4922 : AO221X1 port map( IN1 => RAM_8_26_port, IN2 => n4557, IN3 => 
                           RAM_9_26_port, IN4 => n4546, IN5 => n3681, Q => 
                           n3688);
   U4923 : AO22X1 port map( IN1 => RAM_15_26_port, IN2 => n4579, IN3 => 
                           RAM_14_26_port, IN4 => n4568, Q => n3682);
   U4924 : AO221X1 port map( IN1 => RAM_12_26_port, IN2 => n4601, IN3 => 
                           RAM_13_26_port, IN4 => n4590, IN5 => n3682, Q => 
                           n3687);
   U4925 : AO22X1 port map( IN1 => RAM_3_26_port, IN2 => n4623, IN3 => 
                           RAM_2_26_port, IN4 => n4612, Q => n3683);
   U4926 : AO221X1 port map( IN1 => RAM_0_26_port, IN2 => n4645, IN3 => 
                           RAM_1_26_port, IN4 => n4634, IN5 => n3683, Q => 
                           n3686);
   U4927 : AO22X1 port map( IN1 => RAM_7_26_port, IN2 => n4667, IN3 => 
                           RAM_6_26_port, IN4 => n4656, Q => n3684);
   U4928 : AO221X1 port map( IN1 => RAM_4_26_port, IN2 => n4689, IN3 => 
                           RAM_5_26_port, IN4 => n4678, IN5 => n3684, Q => 
                           n3685);
   U4929 : OR4X1 port map( IN1 => n3688, IN2 => n3687, IN3 => n3686, IN4 => 
                           n3685, Q => RAMDOUT2(26));
   U4930 : AO22X1 port map( IN1 => RAM_11_27_port, IN2 => n4535, IN3 => 
                           RAM_10_27_port, IN4 => n4524, Q => n3689);
   U4931 : AO221X1 port map( IN1 => RAM_8_27_port, IN2 => n4557, IN3 => 
                           RAM_9_27_port, IN4 => n4546, IN5 => n3689, Q => 
                           n3696);
   U4932 : AO22X1 port map( IN1 => RAM_15_27_port, IN2 => n4579, IN3 => 
                           RAM_14_27_port, IN4 => n4568, Q => n3690);
   U4933 : AO221X1 port map( IN1 => RAM_12_27_port, IN2 => n4601, IN3 => 
                           RAM_13_27_port, IN4 => n4590, IN5 => n3690, Q => 
                           n3695);
   U4934 : AO22X1 port map( IN1 => RAM_3_27_port, IN2 => n4623, IN3 => 
                           RAM_2_27_port, IN4 => n4612, Q => n3691);
   U4935 : AO221X1 port map( IN1 => RAM_0_27_port, IN2 => n4645, IN3 => 
                           RAM_1_27_port, IN4 => n4634, IN5 => n3691, Q => 
                           n3694);
   U4936 : AO22X1 port map( IN1 => RAM_7_27_port, IN2 => n4667, IN3 => 
                           RAM_6_27_port, IN4 => n4656, Q => n3692);
   U4937 : AO221X1 port map( IN1 => RAM_4_27_port, IN2 => n4689, IN3 => 
                           RAM_5_27_port, IN4 => n4678, IN5 => n3692, Q => 
                           n3693);
   U4938 : OR4X1 port map( IN1 => n3696, IN2 => n3695, IN3 => n3694, IN4 => 
                           n3693, Q => RAMDOUT2(27));
   U4939 : AO22X1 port map( IN1 => RAM_11_28_port, IN2 => n4535, IN3 => 
                           RAM_10_28_port, IN4 => n4524, Q => n3697);
   U4940 : AO221X1 port map( IN1 => RAM_8_28_port, IN2 => n4557, IN3 => 
                           RAM_9_28_port, IN4 => n4546, IN5 => n3697, Q => 
                           n3704);
   U4941 : AO22X1 port map( IN1 => RAM_15_28_port, IN2 => n4579, IN3 => 
                           RAM_14_28_port, IN4 => n4568, Q => n3698);
   U4942 : AO221X1 port map( IN1 => RAM_12_28_port, IN2 => n4601, IN3 => 
                           RAM_13_28_port, IN4 => n4590, IN5 => n3698, Q => 
                           n3703);
   U4943 : AO22X1 port map( IN1 => RAM_3_28_port, IN2 => n4623, IN3 => 
                           RAM_2_28_port, IN4 => n4612, Q => n3699);
   U4944 : AO221X1 port map( IN1 => RAM_0_28_port, IN2 => n4645, IN3 => 
                           RAM_1_28_port, IN4 => n4634, IN5 => n3699, Q => 
                           n3702);
   U4945 : AO22X1 port map( IN1 => RAM_7_28_port, IN2 => n4667, IN3 => 
                           RAM_6_28_port, IN4 => n4656, Q => n3700);
   U4946 : AO221X1 port map( IN1 => RAM_4_28_port, IN2 => n4689, IN3 => 
                           RAM_5_28_port, IN4 => n4678, IN5 => n3700, Q => 
                           n3701);
   U4947 : OR4X1 port map( IN1 => n3704, IN2 => n3703, IN3 => n3702, IN4 => 
                           n3701, Q => RAMDOUT2(28));
   U4948 : AO22X1 port map( IN1 => RAM_11_29_port, IN2 => n4535, IN3 => 
                           RAM_10_29_port, IN4 => n4524, Q => n3705);
   U4949 : AO221X1 port map( IN1 => RAM_8_29_port, IN2 => n4557, IN3 => 
                           RAM_9_29_port, IN4 => n4546, IN5 => n3705, Q => 
                           n3712);
   U4950 : AO22X1 port map( IN1 => RAM_15_29_port, IN2 => n4579, IN3 => 
                           RAM_14_29_port, IN4 => n4568, Q => n3706);
   U4951 : AO221X1 port map( IN1 => RAM_12_29_port, IN2 => n4601, IN3 => 
                           RAM_13_29_port, IN4 => n4590, IN5 => n3706, Q => 
                           n3711);
   U4952 : AO22X1 port map( IN1 => RAM_3_29_port, IN2 => n4623, IN3 => 
                           RAM_2_29_port, IN4 => n4612, Q => n3707);
   U4953 : AO221X1 port map( IN1 => RAM_0_29_port, IN2 => n4645, IN3 => 
                           RAM_1_29_port, IN4 => n4634, IN5 => n3707, Q => 
                           n3710);
   U4954 : AO22X1 port map( IN1 => RAM_7_29_port, IN2 => n4667, IN3 => 
                           RAM_6_29_port, IN4 => n4656, Q => n3708);
   U4955 : AO221X1 port map( IN1 => RAM_4_29_port, IN2 => n4689, IN3 => 
                           RAM_5_29_port, IN4 => n4678, IN5 => n3708, Q => 
                           n3709);
   U4956 : OR4X1 port map( IN1 => n3712, IN2 => n3711, IN3 => n3710, IN4 => 
                           n3709, Q => RAMDOUT2(29));
   U4957 : AO22X1 port map( IN1 => RAM_11_30_port, IN2 => n4535, IN3 => 
                           RAM_10_30_port, IN4 => n4524, Q => n3713);
   U4958 : AO221X1 port map( IN1 => RAM_8_30_port, IN2 => n4557, IN3 => 
                           RAM_9_30_port, IN4 => n4546, IN5 => n3713, Q => 
                           n3720);
   U4959 : AO22X1 port map( IN1 => RAM_15_30_port, IN2 => n4579, IN3 => 
                           RAM_14_30_port, IN4 => n4568, Q => n3714);
   U4960 : AO221X1 port map( IN1 => RAM_12_30_port, IN2 => n4601, IN3 => 
                           RAM_13_30_port, IN4 => n4590, IN5 => n3714, Q => 
                           n3719);
   U4961 : AO22X1 port map( IN1 => RAM_3_30_port, IN2 => n4623, IN3 => 
                           RAM_2_30_port, IN4 => n4612, Q => n3715);
   U4962 : AO221X1 port map( IN1 => RAM_0_30_port, IN2 => n4645, IN3 => 
                           RAM_1_30_port, IN4 => n4634, IN5 => n3715, Q => 
                           n3718);
   U4963 : AO22X1 port map( IN1 => RAM_7_30_port, IN2 => n4667, IN3 => 
                           RAM_6_30_port, IN4 => n4656, Q => n3716);
   U4964 : AO221X1 port map( IN1 => RAM_4_30_port, IN2 => n4689, IN3 => 
                           RAM_5_30_port, IN4 => n4678, IN5 => n3716, Q => 
                           n3717);
   U4965 : OR4X1 port map( IN1 => n3720, IN2 => n3719, IN3 => n3718, IN4 => 
                           n3717, Q => RAMDOUT2(30));
   U4966 : AO22X1 port map( IN1 => RAM_11_31_port, IN2 => n4535, IN3 => 
                           RAM_10_31_port, IN4 => n4524, Q => n3721);
   U4967 : AO221X1 port map( IN1 => RAM_8_31_port, IN2 => n4557, IN3 => 
                           RAM_9_31_port, IN4 => n4546, IN5 => n3721, Q => 
                           n3728);
   U4968 : AO22X1 port map( IN1 => RAM_15_31_port, IN2 => n4579, IN3 => 
                           RAM_14_31_port, IN4 => n4568, Q => n3722);
   U4969 : AO221X1 port map( IN1 => RAM_12_31_port, IN2 => n4601, IN3 => 
                           RAM_13_31_port, IN4 => n4590, IN5 => n3722, Q => 
                           n3727);
   U4970 : AO22X1 port map( IN1 => RAM_3_31_port, IN2 => n4623, IN3 => 
                           RAM_2_31_port, IN4 => n4612, Q => n3723);
   U4971 : AO221X1 port map( IN1 => RAM_0_31_port, IN2 => n4645, IN3 => 
                           RAM_1_31_port, IN4 => n4634, IN5 => n3723, Q => 
                           n3726);
   U4972 : AO22X1 port map( IN1 => RAM_7_31_port, IN2 => n4667, IN3 => 
                           RAM_6_31_port, IN4 => n4656, Q => n3724);
   U4973 : AO221X1 port map( IN1 => RAM_4_31_port, IN2 => n4689, IN3 => 
                           RAM_5_31_port, IN4 => n4678, IN5 => n3724, Q => 
                           n3725);
   U4974 : OR4X1 port map( IN1 => n3728, IN2 => n3727, IN3 => n3726, IN4 => 
                           n3725, Q => RAMDOUT2(31));
   U4975 : AO22X1 port map( IN1 => RAM_11_32_port, IN2 => n4535, IN3 => 
                           RAM_10_32_port, IN4 => n4524, Q => n3729);
   U4976 : AO221X1 port map( IN1 => RAM_8_32_port, IN2 => n4557, IN3 => 
                           RAM_9_32_port, IN4 => n4546, IN5 => n3729, Q => 
                           n3736);
   U4977 : AO22X1 port map( IN1 => RAM_15_32_port, IN2 => n4579, IN3 => 
                           RAM_14_32_port, IN4 => n4568, Q => n3730);
   U4978 : AO221X1 port map( IN1 => RAM_12_32_port, IN2 => n4601, IN3 => 
                           RAM_13_32_port, IN4 => n4590, IN5 => n3730, Q => 
                           n3735);
   U4979 : AO22X1 port map( IN1 => RAM_3_32_port, IN2 => n4623, IN3 => 
                           RAM_2_32_port, IN4 => n4612, Q => n3731);
   U4980 : AO221X1 port map( IN1 => RAM_0_32_port, IN2 => n4645, IN3 => 
                           RAM_1_32_port, IN4 => n4634, IN5 => n3731, Q => 
                           n3734);
   U4981 : AO22X1 port map( IN1 => RAM_7_32_port, IN2 => n4667, IN3 => 
                           RAM_6_32_port, IN4 => n4656, Q => n3732);
   U4982 : AO221X1 port map( IN1 => RAM_4_32_port, IN2 => n4689, IN3 => 
                           RAM_5_32_port, IN4 => n4678, IN5 => n3732, Q => 
                           n3733);
   U4983 : OR4X1 port map( IN1 => n3736, IN2 => n3735, IN3 => n3734, IN4 => 
                           n3733, Q => RAMDOUT2(32));
   U4984 : AO22X1 port map( IN1 => RAM_11_33_port, IN2 => n4535, IN3 => 
                           RAM_10_33_port, IN4 => n4524, Q => n3737);
   U4985 : AO221X1 port map( IN1 => RAM_8_33_port, IN2 => n4557, IN3 => 
                           RAM_9_33_port, IN4 => n4546, IN5 => n3737, Q => 
                           n3744);
   U4986 : AO22X1 port map( IN1 => RAM_15_33_port, IN2 => n4579, IN3 => 
                           RAM_14_33_port, IN4 => n4568, Q => n3738);
   U4987 : AO221X1 port map( IN1 => RAM_12_33_port, IN2 => n4601, IN3 => 
                           RAM_13_33_port, IN4 => n4590, IN5 => n3738, Q => 
                           n3743);
   U4988 : AO22X1 port map( IN1 => RAM_3_33_port, IN2 => n4623, IN3 => 
                           RAM_2_33_port, IN4 => n4612, Q => n3739);
   U4989 : AO221X1 port map( IN1 => RAM_0_33_port, IN2 => n4645, IN3 => 
                           RAM_1_33_port, IN4 => n4634, IN5 => n3739, Q => 
                           n3742);
   U4990 : AO22X1 port map( IN1 => RAM_7_33_port, IN2 => n4667, IN3 => 
                           RAM_6_33_port, IN4 => n4656, Q => n3740);
   U4991 : AO221X1 port map( IN1 => RAM_4_33_port, IN2 => n4689, IN3 => 
                           RAM_5_33_port, IN4 => n4678, IN5 => n3740, Q => 
                           n3741);
   U4992 : OR4X1 port map( IN1 => n3744, IN2 => n3743, IN3 => n3742, IN4 => 
                           n3741, Q => RAMDOUT2(33));
   U4993 : AO22X1 port map( IN1 => RAM_11_34_port, IN2 => n4535, IN3 => 
                           RAM_10_34_port, IN4 => n4524, Q => n3745);
   U4994 : AO221X1 port map( IN1 => RAM_8_34_port, IN2 => n4557, IN3 => 
                           RAM_9_34_port, IN4 => n4546, IN5 => n3745, Q => 
                           n3752);
   U4995 : AO22X1 port map( IN1 => RAM_15_34_port, IN2 => n4579, IN3 => 
                           RAM_14_34_port, IN4 => n4568, Q => n3746);
   U4996 : AO221X1 port map( IN1 => RAM_12_34_port, IN2 => n4601, IN3 => 
                           RAM_13_34_port, IN4 => n4590, IN5 => n3746, Q => 
                           n3751);
   U4997 : AO22X1 port map( IN1 => RAM_3_34_port, IN2 => n4623, IN3 => 
                           RAM_2_34_port, IN4 => n4612, Q => n3747);
   U4998 : AO221X1 port map( IN1 => RAM_0_34_port, IN2 => n4645, IN3 => 
                           RAM_1_34_port, IN4 => n4634, IN5 => n3747, Q => 
                           n3750);
   U4999 : AO22X1 port map( IN1 => RAM_7_34_port, IN2 => n4667, IN3 => 
                           RAM_6_34_port, IN4 => n4656, Q => n3748);
   U5000 : AO221X1 port map( IN1 => RAM_4_34_port, IN2 => n4689, IN3 => 
                           RAM_5_34_port, IN4 => n4678, IN5 => n3748, Q => 
                           n3749);
   U5001 : OR4X1 port map( IN1 => n3752, IN2 => n3751, IN3 => n3750, IN4 => 
                           n3749, Q => RAMDOUT2(34));
   U5002 : AO22X1 port map( IN1 => RAM_11_35_port, IN2 => n4535, IN3 => 
                           RAM_10_35_port, IN4 => n4524, Q => n3753);
   U5003 : AO221X1 port map( IN1 => RAM_8_35_port, IN2 => n4557, IN3 => 
                           RAM_9_35_port, IN4 => n4546, IN5 => n3753, Q => 
                           n3760);
   U5004 : AO22X1 port map( IN1 => RAM_15_35_port, IN2 => n4579, IN3 => 
                           RAM_14_35_port, IN4 => n4568, Q => n3754);
   U5005 : AO221X1 port map( IN1 => RAM_12_35_port, IN2 => n4601, IN3 => 
                           RAM_13_35_port, IN4 => n4590, IN5 => n3754, Q => 
                           n3759);
   U5006 : AO22X1 port map( IN1 => RAM_3_35_port, IN2 => n4623, IN3 => 
                           RAM_2_35_port, IN4 => n4612, Q => n3755);
   U5007 : AO221X1 port map( IN1 => RAM_0_35_port, IN2 => n4645, IN3 => 
                           RAM_1_35_port, IN4 => n4634, IN5 => n3755, Q => 
                           n3758);
   U5008 : AO22X1 port map( IN1 => RAM_7_35_port, IN2 => n4667, IN3 => 
                           RAM_6_35_port, IN4 => n4656, Q => n3756);
   U5009 : AO221X1 port map( IN1 => RAM_4_35_port, IN2 => n4689, IN3 => 
                           RAM_5_35_port, IN4 => n4678, IN5 => n3756, Q => 
                           n3757);
   U5010 : OR4X1 port map( IN1 => n3760, IN2 => n3759, IN3 => n3758, IN4 => 
                           n3757, Q => RAMDOUT2(35));
   U5011 : AO22X1 port map( IN1 => RAM_11_36_port, IN2 => n4534, IN3 => 
                           RAM_10_36_port, IN4 => n4523, Q => n3761);
   U5012 : AO221X1 port map( IN1 => RAM_8_36_port, IN2 => n4556, IN3 => 
                           RAM_9_36_port, IN4 => n4545, IN5 => n3761, Q => 
                           n3768);
   U5013 : AO22X1 port map( IN1 => RAM_15_36_port, IN2 => n4578, IN3 => 
                           RAM_14_36_port, IN4 => n4567, Q => n3762);
   U5014 : AO221X1 port map( IN1 => RAM_12_36_port, IN2 => n4600, IN3 => 
                           RAM_13_36_port, IN4 => n4589, IN5 => n3762, Q => 
                           n3767);
   U5015 : AO22X1 port map( IN1 => RAM_3_36_port, IN2 => n4622, IN3 => 
                           RAM_2_36_port, IN4 => n4611, Q => n3763);
   U5016 : AO221X1 port map( IN1 => RAM_0_36_port, IN2 => n4644, IN3 => 
                           RAM_1_36_port, IN4 => n4633, IN5 => n3763, Q => 
                           n3766);
   U5017 : AO22X1 port map( IN1 => RAM_7_36_port, IN2 => n4666, IN3 => 
                           RAM_6_36_port, IN4 => n4655, Q => n3764);
   U5018 : AO221X1 port map( IN1 => RAM_4_36_port, IN2 => n4688, IN3 => 
                           RAM_5_36_port, IN4 => n4677, IN5 => n3764, Q => 
                           n3765);
   U5019 : OR4X1 port map( IN1 => n3768, IN2 => n3767, IN3 => n3766, IN4 => 
                           n3765, Q => RAMDOUT2(36));
   U5020 : AO22X1 port map( IN1 => RAM_11_37_port, IN2 => n4534, IN3 => 
                           RAM_10_37_port, IN4 => n4523, Q => n3769);
   U5021 : AO221X1 port map( IN1 => RAM_8_37_port, IN2 => n4556, IN3 => 
                           RAM_9_37_port, IN4 => n4545, IN5 => n3769, Q => 
                           n3776);
   U5022 : AO22X1 port map( IN1 => RAM_15_37_port, IN2 => n4578, IN3 => 
                           RAM_14_37_port, IN4 => n4567, Q => n3770);
   U5023 : AO221X1 port map( IN1 => RAM_12_37_port, IN2 => n4600, IN3 => 
                           RAM_13_37_port, IN4 => n4589, IN5 => n3770, Q => 
                           n3775);
   U5024 : AO22X1 port map( IN1 => RAM_3_37_port, IN2 => n4622, IN3 => 
                           RAM_2_37_port, IN4 => n4611, Q => n3771);
   U5025 : AO221X1 port map( IN1 => RAM_0_37_port, IN2 => n4644, IN3 => 
                           RAM_1_37_port, IN4 => n4633, IN5 => n3771, Q => 
                           n3774);
   U5026 : AO22X1 port map( IN1 => RAM_7_37_port, IN2 => n4666, IN3 => 
                           RAM_6_37_port, IN4 => n4655, Q => n3772);
   U5027 : AO221X1 port map( IN1 => RAM_4_37_port, IN2 => n4688, IN3 => 
                           RAM_5_37_port, IN4 => n4677, IN5 => n3772, Q => 
                           n3773);
   U5028 : OR4X1 port map( IN1 => n3776, IN2 => n3775, IN3 => n3774, IN4 => 
                           n3773, Q => RAMDOUT2(37));
   U5029 : AO22X1 port map( IN1 => RAM_11_38_port, IN2 => n4534, IN3 => 
                           RAM_10_38_port, IN4 => n4523, Q => n3777);
   U5030 : AO221X1 port map( IN1 => RAM_8_38_port, IN2 => n4556, IN3 => 
                           RAM_9_38_port, IN4 => n4545, IN5 => n3777, Q => 
                           n3784);
   U5031 : AO22X1 port map( IN1 => RAM_15_38_port, IN2 => n4578, IN3 => 
                           RAM_14_38_port, IN4 => n4567, Q => n3778);
   U5032 : AO221X1 port map( IN1 => RAM_12_38_port, IN2 => n4600, IN3 => 
                           RAM_13_38_port, IN4 => n4589, IN5 => n3778, Q => 
                           n3783);
   U5033 : AO22X1 port map( IN1 => RAM_3_38_port, IN2 => n4622, IN3 => 
                           RAM_2_38_port, IN4 => n4611, Q => n3779);
   U5034 : AO221X1 port map( IN1 => RAM_0_38_port, IN2 => n4644, IN3 => 
                           RAM_1_38_port, IN4 => n4633, IN5 => n3779, Q => 
                           n3782);
   U5035 : AO22X1 port map( IN1 => RAM_7_38_port, IN2 => n4666, IN3 => 
                           RAM_6_38_port, IN4 => n4655, Q => n3780);
   U5036 : AO221X1 port map( IN1 => RAM_4_38_port, IN2 => n4688, IN3 => 
                           RAM_5_38_port, IN4 => n4677, IN5 => n3780, Q => 
                           n3781);
   U5037 : OR4X1 port map( IN1 => n3784, IN2 => n3783, IN3 => n3782, IN4 => 
                           n3781, Q => RAMDOUT2(38));
   U5038 : AO22X1 port map( IN1 => RAM_11_39_port, IN2 => n4534, IN3 => 
                           RAM_10_39_port, IN4 => n4523, Q => n3785);
   U5039 : AO221X1 port map( IN1 => RAM_8_39_port, IN2 => n4556, IN3 => 
                           RAM_9_39_port, IN4 => n4545, IN5 => n3785, Q => 
                           n3792);
   U5040 : AO22X1 port map( IN1 => RAM_15_39_port, IN2 => n4578, IN3 => 
                           RAM_14_39_port, IN4 => n4567, Q => n3786);
   U5041 : AO221X1 port map( IN1 => RAM_12_39_port, IN2 => n4600, IN3 => 
                           RAM_13_39_port, IN4 => n4589, IN5 => n3786, Q => 
                           n3791);
   U5042 : AO22X1 port map( IN1 => RAM_3_39_port, IN2 => n4622, IN3 => 
                           RAM_2_39_port, IN4 => n4611, Q => n3787);
   U5043 : AO221X1 port map( IN1 => RAM_0_39_port, IN2 => n4644, IN3 => 
                           RAM_1_39_port, IN4 => n4633, IN5 => n3787, Q => 
                           n3790);
   U5044 : AO22X1 port map( IN1 => RAM_7_39_port, IN2 => n4666, IN3 => 
                           RAM_6_39_port, IN4 => n4655, Q => n3788);
   U5045 : AO221X1 port map( IN1 => RAM_4_39_port, IN2 => n4688, IN3 => 
                           RAM_5_39_port, IN4 => n4677, IN5 => n3788, Q => 
                           n3789);
   U5046 : OR4X1 port map( IN1 => n3792, IN2 => n3791, IN3 => n3790, IN4 => 
                           n3789, Q => RAMDOUT2(39));
   U5047 : AO22X1 port map( IN1 => RAM_11_40_port, IN2 => n4534, IN3 => 
                           RAM_10_40_port, IN4 => n4523, Q => n3793);
   U5048 : AO221X1 port map( IN1 => RAM_8_40_port, IN2 => n4556, IN3 => 
                           RAM_9_40_port, IN4 => n4545, IN5 => n3793, Q => 
                           n3800);
   U5049 : AO22X1 port map( IN1 => RAM_15_40_port, IN2 => n4578, IN3 => 
                           RAM_14_40_port, IN4 => n4567, Q => n3794);
   U5050 : AO221X1 port map( IN1 => RAM_12_40_port, IN2 => n4600, IN3 => 
                           RAM_13_40_port, IN4 => n4589, IN5 => n3794, Q => 
                           n3799);
   U5051 : AO22X1 port map( IN1 => RAM_3_40_port, IN2 => n4622, IN3 => 
                           RAM_2_40_port, IN4 => n4611, Q => n3795);
   U5052 : AO221X1 port map( IN1 => RAM_0_40_port, IN2 => n4644, IN3 => 
                           RAM_1_40_port, IN4 => n4633, IN5 => n3795, Q => 
                           n3798);
   U5053 : AO22X1 port map( IN1 => RAM_7_40_port, IN2 => n4666, IN3 => 
                           RAM_6_40_port, IN4 => n4655, Q => n3796);
   U5054 : AO221X1 port map( IN1 => RAM_4_40_port, IN2 => n4688, IN3 => 
                           RAM_5_40_port, IN4 => n4677, IN5 => n3796, Q => 
                           n3797);
   U5055 : OR4X1 port map( IN1 => n3800, IN2 => n3799, IN3 => n3798, IN4 => 
                           n3797, Q => RAMDOUT2(40));
   U5056 : AO22X1 port map( IN1 => RAM_11_41_port, IN2 => n4534, IN3 => 
                           RAM_10_41_port, IN4 => n4523, Q => n3801);
   U5057 : AO221X1 port map( IN1 => RAM_8_41_port, IN2 => n4556, IN3 => 
                           RAM_9_41_port, IN4 => n4545, IN5 => n3801, Q => 
                           n3808);
   U5058 : AO22X1 port map( IN1 => RAM_15_41_port, IN2 => n4578, IN3 => 
                           RAM_14_41_port, IN4 => n4567, Q => n3802);
   U5059 : AO221X1 port map( IN1 => RAM_12_41_port, IN2 => n4600, IN3 => 
                           RAM_13_41_port, IN4 => n4589, IN5 => n3802, Q => 
                           n3807);
   U5060 : AO22X1 port map( IN1 => RAM_3_41_port, IN2 => n4622, IN3 => 
                           RAM_2_41_port, IN4 => n4611, Q => n3803);
   U5061 : AO221X1 port map( IN1 => RAM_0_41_port, IN2 => n4644, IN3 => 
                           RAM_1_41_port, IN4 => n4633, IN5 => n3803, Q => 
                           n3806);
   U5062 : AO22X1 port map( IN1 => RAM_7_41_port, IN2 => n4666, IN3 => 
                           RAM_6_41_port, IN4 => n4655, Q => n3804);
   U5063 : AO221X1 port map( IN1 => RAM_4_41_port, IN2 => n4688, IN3 => 
                           RAM_5_41_port, IN4 => n4677, IN5 => n3804, Q => 
                           n3805);
   U5064 : OR4X1 port map( IN1 => n3808, IN2 => n3807, IN3 => n3806, IN4 => 
                           n3805, Q => RAMDOUT2(41));
   U5065 : AO22X1 port map( IN1 => RAM_11_42_port, IN2 => n4534, IN3 => 
                           RAM_10_42_port, IN4 => n4523, Q => n3809);
   U5066 : AO221X1 port map( IN1 => RAM_8_42_port, IN2 => n4556, IN3 => 
                           RAM_9_42_port, IN4 => n4545, IN5 => n3809, Q => 
                           n3816);
   U5067 : AO22X1 port map( IN1 => RAM_15_42_port, IN2 => n4578, IN3 => 
                           RAM_14_42_port, IN4 => n4567, Q => n3810);
   U5068 : AO221X1 port map( IN1 => RAM_12_42_port, IN2 => n4600, IN3 => 
                           RAM_13_42_port, IN4 => n4589, IN5 => n3810, Q => 
                           n3815);
   U5069 : AO22X1 port map( IN1 => RAM_3_42_port, IN2 => n4622, IN3 => 
                           RAM_2_42_port, IN4 => n4611, Q => n3811);
   U5070 : AO221X1 port map( IN1 => RAM_0_42_port, IN2 => n4644, IN3 => 
                           RAM_1_42_port, IN4 => n4633, IN5 => n3811, Q => 
                           n3814);
   U5071 : AO22X1 port map( IN1 => RAM_7_42_port, IN2 => n4666, IN3 => 
                           RAM_6_42_port, IN4 => n4655, Q => n3812);
   U5072 : AO221X1 port map( IN1 => RAM_4_42_port, IN2 => n4688, IN3 => 
                           RAM_5_42_port, IN4 => n4677, IN5 => n3812, Q => 
                           n3813);
   U5073 : OR4X1 port map( IN1 => n3816, IN2 => n3815, IN3 => n3814, IN4 => 
                           n3813, Q => RAMDOUT2(42));
   U5074 : AO22X1 port map( IN1 => RAM_11_43_port, IN2 => n4534, IN3 => 
                           RAM_10_43_port, IN4 => n4523, Q => n3817);
   U5075 : AO221X1 port map( IN1 => RAM_8_43_port, IN2 => n4556, IN3 => 
                           RAM_9_43_port, IN4 => n4545, IN5 => n3817, Q => 
                           n3824);
   U5076 : AO22X1 port map( IN1 => RAM_15_43_port, IN2 => n4578, IN3 => 
                           RAM_14_43_port, IN4 => n4567, Q => n3818);
   U5077 : AO221X1 port map( IN1 => RAM_12_43_port, IN2 => n4600, IN3 => 
                           RAM_13_43_port, IN4 => n4589, IN5 => n3818, Q => 
                           n3823);
   U5078 : AO22X1 port map( IN1 => RAM_3_43_port, IN2 => n4622, IN3 => 
                           RAM_2_43_port, IN4 => n4611, Q => n3819);
   U5079 : AO221X1 port map( IN1 => RAM_0_43_port, IN2 => n4644, IN3 => 
                           RAM_1_43_port, IN4 => n4633, IN5 => n3819, Q => 
                           n3822);
   U5080 : AO22X1 port map( IN1 => RAM_7_43_port, IN2 => n4666, IN3 => 
                           RAM_6_43_port, IN4 => n4655, Q => n3820);
   U5081 : AO221X1 port map( IN1 => RAM_4_43_port, IN2 => n4688, IN3 => 
                           RAM_5_43_port, IN4 => n4677, IN5 => n3820, Q => 
                           n3821);
   U5082 : OR4X1 port map( IN1 => n3824, IN2 => n3823, IN3 => n3822, IN4 => 
                           n3821, Q => RAMDOUT2(43));
   U5083 : AO22X1 port map( IN1 => RAM_11_44_port, IN2 => n4534, IN3 => 
                           RAM_10_44_port, IN4 => n4523, Q => n3825);
   U5084 : AO221X1 port map( IN1 => RAM_8_44_port, IN2 => n4556, IN3 => 
                           RAM_9_44_port, IN4 => n4545, IN5 => n3825, Q => 
                           n3832);
   U5085 : AO22X1 port map( IN1 => RAM_15_44_port, IN2 => n4578, IN3 => 
                           RAM_14_44_port, IN4 => n4567, Q => n3826);
   U5086 : AO221X1 port map( IN1 => RAM_12_44_port, IN2 => n4600, IN3 => 
                           RAM_13_44_port, IN4 => n4589, IN5 => n3826, Q => 
                           n3831);
   U5087 : AO22X1 port map( IN1 => RAM_3_44_port, IN2 => n4622, IN3 => 
                           RAM_2_44_port, IN4 => n4611, Q => n3827);
   U5088 : AO221X1 port map( IN1 => RAM_0_44_port, IN2 => n4644, IN3 => 
                           RAM_1_44_port, IN4 => n4633, IN5 => n3827, Q => 
                           n3830);
   U5089 : AO22X1 port map( IN1 => RAM_7_44_port, IN2 => n4666, IN3 => 
                           RAM_6_44_port, IN4 => n4655, Q => n3828);
   U5090 : AO221X1 port map( IN1 => RAM_4_44_port, IN2 => n4688, IN3 => 
                           RAM_5_44_port, IN4 => n4677, IN5 => n3828, Q => 
                           n3829);
   U5091 : OR4X1 port map( IN1 => n3832, IN2 => n3831, IN3 => n3830, IN4 => 
                           n3829, Q => RAMDOUT2(44));
   U5092 : AO22X1 port map( IN1 => RAM_11_45_port, IN2 => n4534, IN3 => 
                           RAM_10_45_port, IN4 => n4523, Q => n3833);
   U5093 : AO221X1 port map( IN1 => RAM_8_45_port, IN2 => n4556, IN3 => 
                           RAM_9_45_port, IN4 => n4545, IN5 => n3833, Q => 
                           n3840);
   U5094 : AO22X1 port map( IN1 => RAM_15_45_port, IN2 => n4578, IN3 => 
                           RAM_14_45_port, IN4 => n4567, Q => n3834);
   U5095 : AO221X1 port map( IN1 => RAM_12_45_port, IN2 => n4600, IN3 => 
                           RAM_13_45_port, IN4 => n4589, IN5 => n3834, Q => 
                           n3839);
   U5096 : AO22X1 port map( IN1 => RAM_3_45_port, IN2 => n4622, IN3 => 
                           RAM_2_45_port, IN4 => n4611, Q => n3835);
   U5097 : AO221X1 port map( IN1 => RAM_0_45_port, IN2 => n4644, IN3 => 
                           RAM_1_45_port, IN4 => n4633, IN5 => n3835, Q => 
                           n3838);
   U5098 : AO22X1 port map( IN1 => RAM_7_45_port, IN2 => n4666, IN3 => 
                           RAM_6_45_port, IN4 => n4655, Q => n3836);
   U5099 : AO221X1 port map( IN1 => RAM_4_45_port, IN2 => n4688, IN3 => 
                           RAM_5_45_port, IN4 => n4677, IN5 => n3836, Q => 
                           n3837);
   U5100 : OR4X1 port map( IN1 => n3840, IN2 => n3839, IN3 => n3838, IN4 => 
                           n3837, Q => RAMDOUT2(45));
   U5101 : AO22X1 port map( IN1 => RAM_11_46_port, IN2 => n4534, IN3 => 
                           RAM_10_46_port, IN4 => n4523, Q => n3841);
   U5102 : AO221X1 port map( IN1 => RAM_8_46_port, IN2 => n4556, IN3 => 
                           RAM_9_46_port, IN4 => n4545, IN5 => n3841, Q => 
                           n3848);
   U5103 : AO22X1 port map( IN1 => RAM_15_46_port, IN2 => n4578, IN3 => 
                           RAM_14_46_port, IN4 => n4567, Q => n3842);
   U5104 : AO221X1 port map( IN1 => RAM_12_46_port, IN2 => n4600, IN3 => 
                           RAM_13_46_port, IN4 => n4589, IN5 => n3842, Q => 
                           n3847);
   U5105 : AO22X1 port map( IN1 => RAM_3_46_port, IN2 => n4622, IN3 => 
                           RAM_2_46_port, IN4 => n4611, Q => n3843);
   U5106 : AO221X1 port map( IN1 => RAM_0_46_port, IN2 => n4644, IN3 => 
                           RAM_1_46_port, IN4 => n4633, IN5 => n3843, Q => 
                           n3846);
   U5107 : AO22X1 port map( IN1 => RAM_7_46_port, IN2 => n4666, IN3 => 
                           RAM_6_46_port, IN4 => n4655, Q => n3844);
   U5108 : AO221X1 port map( IN1 => RAM_4_46_port, IN2 => n4688, IN3 => 
                           RAM_5_46_port, IN4 => n4677, IN5 => n3844, Q => 
                           n3845);
   U5109 : OR4X1 port map( IN1 => n3848, IN2 => n3847, IN3 => n3846, IN4 => 
                           n3845, Q => RAMDOUT2(46));
   U5110 : AO22X1 port map( IN1 => RAM_11_47_port, IN2 => n4534, IN3 => 
                           RAM_10_47_port, IN4 => n4523, Q => n3849);
   U5111 : AO221X1 port map( IN1 => RAM_8_47_port, IN2 => n4556, IN3 => 
                           RAM_9_47_port, IN4 => n4545, IN5 => n3849, Q => 
                           n3856);
   U5112 : AO22X1 port map( IN1 => RAM_15_47_port, IN2 => n4578, IN3 => 
                           RAM_14_47_port, IN4 => n4567, Q => n3850);
   U5113 : AO221X1 port map( IN1 => RAM_12_47_port, IN2 => n4600, IN3 => 
                           RAM_13_47_port, IN4 => n4589, IN5 => n3850, Q => 
                           n3855);
   U5114 : AO22X1 port map( IN1 => RAM_3_47_port, IN2 => n4622, IN3 => 
                           RAM_2_47_port, IN4 => n4611, Q => n3851);
   U5115 : AO221X1 port map( IN1 => RAM_0_47_port, IN2 => n4644, IN3 => 
                           RAM_1_47_port, IN4 => n4633, IN5 => n3851, Q => 
                           n3854);
   U5116 : AO22X1 port map( IN1 => RAM_7_47_port, IN2 => n4666, IN3 => 
                           RAM_6_47_port, IN4 => n4655, Q => n3852);
   U5117 : AO221X1 port map( IN1 => RAM_4_47_port, IN2 => n4688, IN3 => 
                           RAM_5_47_port, IN4 => n4677, IN5 => n3852, Q => 
                           n3853);
   U5118 : OR4X1 port map( IN1 => n3856, IN2 => n3855, IN3 => n3854, IN4 => 
                           n3853, Q => RAMDOUT2(47));
   U5119 : AO22X1 port map( IN1 => RAM_11_48_port, IN2 => n4533, IN3 => 
                           RAM_10_48_port, IN4 => n4522, Q => n3857);
   U5120 : AO221X1 port map( IN1 => RAM_8_48_port, IN2 => n4555, IN3 => 
                           RAM_9_48_port, IN4 => n4544, IN5 => n3857, Q => 
                           n3864);
   U5121 : AO22X1 port map( IN1 => RAM_15_48_port, IN2 => n4577, IN3 => 
                           RAM_14_48_port, IN4 => n4566, Q => n3858);
   U5122 : AO221X1 port map( IN1 => RAM_12_48_port, IN2 => n4599, IN3 => 
                           RAM_13_48_port, IN4 => n4588, IN5 => n3858, Q => 
                           n3863);
   U5123 : AO22X1 port map( IN1 => RAM_3_48_port, IN2 => n4621, IN3 => 
                           RAM_2_48_port, IN4 => n4610, Q => n3859);
   U5124 : AO221X1 port map( IN1 => RAM_0_48_port, IN2 => n4643, IN3 => 
                           RAM_1_48_port, IN4 => n4632, IN5 => n3859, Q => 
                           n3862);
   U5125 : AO22X1 port map( IN1 => RAM_7_48_port, IN2 => n4665, IN3 => 
                           RAM_6_48_port, IN4 => n4654, Q => n3860);
   U5126 : AO221X1 port map( IN1 => RAM_4_48_port, IN2 => n4687, IN3 => 
                           RAM_5_48_port, IN4 => n4676, IN5 => n3860, Q => 
                           n3861);
   U5127 : OR4X1 port map( IN1 => n3864, IN2 => n3863, IN3 => n3862, IN4 => 
                           n3861, Q => RAMDOUT2(48));
   U5128 : AO22X1 port map( IN1 => RAM_11_49_port, IN2 => n4533, IN3 => 
                           RAM_10_49_port, IN4 => n4522, Q => n3865);
   U5129 : AO221X1 port map( IN1 => RAM_8_49_port, IN2 => n4555, IN3 => 
                           RAM_9_49_port, IN4 => n4544, IN5 => n3865, Q => 
                           n3872);
   U5130 : AO22X1 port map( IN1 => RAM_15_49_port, IN2 => n4577, IN3 => 
                           RAM_14_49_port, IN4 => n4566, Q => n3866);
   U5131 : AO221X1 port map( IN1 => RAM_12_49_port, IN2 => n4599, IN3 => 
                           RAM_13_49_port, IN4 => n4588, IN5 => n3866, Q => 
                           n3871);
   U5132 : AO22X1 port map( IN1 => RAM_3_49_port, IN2 => n4621, IN3 => 
                           RAM_2_49_port, IN4 => n4610, Q => n3867);
   U5133 : AO221X1 port map( IN1 => RAM_0_49_port, IN2 => n4643, IN3 => 
                           RAM_1_49_port, IN4 => n4632, IN5 => n3867, Q => 
                           n3870);
   U5134 : AO22X1 port map( IN1 => RAM_7_49_port, IN2 => n4665, IN3 => 
                           RAM_6_49_port, IN4 => n4654, Q => n3868);
   U5135 : AO221X1 port map( IN1 => RAM_4_49_port, IN2 => n4687, IN3 => 
                           RAM_5_49_port, IN4 => n4676, IN5 => n3868, Q => 
                           n3869);
   U5136 : OR4X1 port map( IN1 => n3872, IN2 => n3871, IN3 => n3870, IN4 => 
                           n3869, Q => RAMDOUT2(49));
   U5137 : AO22X1 port map( IN1 => RAM_11_50_port, IN2 => n4533, IN3 => 
                           RAM_10_50_port, IN4 => n4522, Q => n3873);
   U5138 : AO221X1 port map( IN1 => RAM_8_50_port, IN2 => n4555, IN3 => 
                           RAM_9_50_port, IN4 => n4544, IN5 => n3873, Q => 
                           n3880);
   U5139 : AO22X1 port map( IN1 => RAM_15_50_port, IN2 => n4577, IN3 => 
                           RAM_14_50_port, IN4 => n4566, Q => n3874);
   U5140 : AO221X1 port map( IN1 => RAM_12_50_port, IN2 => n4599, IN3 => 
                           RAM_13_50_port, IN4 => n4588, IN5 => n3874, Q => 
                           n3879);
   U5141 : AO22X1 port map( IN1 => RAM_3_50_port, IN2 => n4621, IN3 => 
                           RAM_2_50_port, IN4 => n4610, Q => n3875);
   U5142 : AO221X1 port map( IN1 => RAM_0_50_port, IN2 => n4643, IN3 => 
                           RAM_1_50_port, IN4 => n4632, IN5 => n3875, Q => 
                           n3878);
   U5143 : AO22X1 port map( IN1 => RAM_7_50_port, IN2 => n4665, IN3 => 
                           RAM_6_50_port, IN4 => n4654, Q => n3876);
   U5144 : AO221X1 port map( IN1 => RAM_4_50_port, IN2 => n4687, IN3 => 
                           RAM_5_50_port, IN4 => n4676, IN5 => n3876, Q => 
                           n3877);
   U5145 : OR4X1 port map( IN1 => n3880, IN2 => n3879, IN3 => n3878, IN4 => 
                           n3877, Q => RAMDOUT2(50));
   U5146 : AO22X1 port map( IN1 => RAM_11_51_port, IN2 => n4533, IN3 => 
                           RAM_10_51_port, IN4 => n4522, Q => n3881);
   U5147 : AO221X1 port map( IN1 => RAM_8_51_port, IN2 => n4555, IN3 => 
                           RAM_9_51_port, IN4 => n4544, IN5 => n3881, Q => 
                           n3888);
   U5148 : AO22X1 port map( IN1 => RAM_15_51_port, IN2 => n4577, IN3 => 
                           RAM_14_51_port, IN4 => n4566, Q => n3882);
   U5149 : AO221X1 port map( IN1 => RAM_12_51_port, IN2 => n4599, IN3 => 
                           RAM_13_51_port, IN4 => n4588, IN5 => n3882, Q => 
                           n3887);
   U5150 : AO22X1 port map( IN1 => RAM_3_51_port, IN2 => n4621, IN3 => 
                           RAM_2_51_port, IN4 => n4610, Q => n3883);
   U5151 : AO221X1 port map( IN1 => RAM_0_51_port, IN2 => n4643, IN3 => 
                           RAM_1_51_port, IN4 => n4632, IN5 => n3883, Q => 
                           n3886);
   U5152 : AO22X1 port map( IN1 => RAM_7_51_port, IN2 => n4665, IN3 => 
                           RAM_6_51_port, IN4 => n4654, Q => n3884);
   U5153 : AO221X1 port map( IN1 => RAM_4_51_port, IN2 => n4687, IN3 => 
                           RAM_5_51_port, IN4 => n4676, IN5 => n3884, Q => 
                           n3885);
   U5154 : OR4X1 port map( IN1 => n3888, IN2 => n3887, IN3 => n3886, IN4 => 
                           n3885, Q => RAMDOUT2(51));
   U5155 : AO22X1 port map( IN1 => RAM_11_52_port, IN2 => n4533, IN3 => 
                           RAM_10_52_port, IN4 => n4522, Q => n3889);
   U5156 : AO221X1 port map( IN1 => RAM_8_52_port, IN2 => n4555, IN3 => 
                           RAM_9_52_port, IN4 => n4544, IN5 => n3889, Q => 
                           n3896);
   U5157 : AO22X1 port map( IN1 => RAM_15_52_port, IN2 => n4577, IN3 => 
                           RAM_14_52_port, IN4 => n4566, Q => n3890);
   U5158 : AO221X1 port map( IN1 => RAM_12_52_port, IN2 => n4599, IN3 => 
                           RAM_13_52_port, IN4 => n4588, IN5 => n3890, Q => 
                           n3895);
   U5159 : AO22X1 port map( IN1 => RAM_3_52_port, IN2 => n4621, IN3 => 
                           RAM_2_52_port, IN4 => n4610, Q => n3891);
   U5160 : AO221X1 port map( IN1 => RAM_0_52_port, IN2 => n4643, IN3 => 
                           RAM_1_52_port, IN4 => n4632, IN5 => n3891, Q => 
                           n3894);
   U5161 : AO22X1 port map( IN1 => RAM_7_52_port, IN2 => n4665, IN3 => 
                           RAM_6_52_port, IN4 => n4654, Q => n3892);
   U5162 : AO221X1 port map( IN1 => RAM_4_52_port, IN2 => n4687, IN3 => 
                           RAM_5_52_port, IN4 => n4676, IN5 => n3892, Q => 
                           n3893);
   U5163 : OR4X1 port map( IN1 => n3896, IN2 => n3895, IN3 => n3894, IN4 => 
                           n3893, Q => RAMDOUT2(52));
   U5164 : AO22X1 port map( IN1 => RAM_11_53_port, IN2 => n4533, IN3 => 
                           RAM_10_53_port, IN4 => n4522, Q => n3897);
   U5165 : AO221X1 port map( IN1 => RAM_8_53_port, IN2 => n4555, IN3 => 
                           RAM_9_53_port, IN4 => n4544, IN5 => n3897, Q => 
                           n3904);
   U5166 : AO22X1 port map( IN1 => RAM_15_53_port, IN2 => n4577, IN3 => 
                           RAM_14_53_port, IN4 => n4566, Q => n3898);
   U5167 : AO221X1 port map( IN1 => RAM_12_53_port, IN2 => n4599, IN3 => 
                           RAM_13_53_port, IN4 => n4588, IN5 => n3898, Q => 
                           n3903);
   U5168 : AO22X1 port map( IN1 => RAM_3_53_port, IN2 => n4621, IN3 => 
                           RAM_2_53_port, IN4 => n4610, Q => n3899);
   U5169 : AO221X1 port map( IN1 => RAM_0_53_port, IN2 => n4643, IN3 => 
                           RAM_1_53_port, IN4 => n4632, IN5 => n3899, Q => 
                           n3902);
   U5170 : AO22X1 port map( IN1 => RAM_7_53_port, IN2 => n4665, IN3 => 
                           RAM_6_53_port, IN4 => n4654, Q => n3900);
   U5171 : AO221X1 port map( IN1 => RAM_4_53_port, IN2 => n4687, IN3 => 
                           RAM_5_53_port, IN4 => n4676, IN5 => n3900, Q => 
                           n3901);
   U5172 : OR4X1 port map( IN1 => n3904, IN2 => n3903, IN3 => n3902, IN4 => 
                           n3901, Q => RAMDOUT2(53));
   U5173 : AO22X1 port map( IN1 => RAM_11_54_port, IN2 => n4533, IN3 => 
                           RAM_10_54_port, IN4 => n4522, Q => n3905);
   U5174 : AO221X1 port map( IN1 => RAM_8_54_port, IN2 => n4555, IN3 => 
                           RAM_9_54_port, IN4 => n4544, IN5 => n3905, Q => 
                           n3912);
   U5175 : AO22X1 port map( IN1 => RAM_15_54_port, IN2 => n4577, IN3 => 
                           RAM_14_54_port, IN4 => n4566, Q => n3906);
   U5176 : AO221X1 port map( IN1 => RAM_12_54_port, IN2 => n4599, IN3 => 
                           RAM_13_54_port, IN4 => n4588, IN5 => n3906, Q => 
                           n3911);
   U5177 : AO22X1 port map( IN1 => RAM_3_54_port, IN2 => n4621, IN3 => 
                           RAM_2_54_port, IN4 => n4610, Q => n3907);
   U5178 : AO221X1 port map( IN1 => RAM_0_54_port, IN2 => n4643, IN3 => 
                           RAM_1_54_port, IN4 => n4632, IN5 => n3907, Q => 
                           n3910);
   U5179 : AO22X1 port map( IN1 => RAM_7_54_port, IN2 => n4665, IN3 => 
                           RAM_6_54_port, IN4 => n4654, Q => n3908);
   U5180 : AO221X1 port map( IN1 => RAM_4_54_port, IN2 => n4687, IN3 => 
                           RAM_5_54_port, IN4 => n4676, IN5 => n3908, Q => 
                           n3909);
   U5181 : OR4X1 port map( IN1 => n3912, IN2 => n3911, IN3 => n3910, IN4 => 
                           n3909, Q => RAMDOUT2(54));
   U5182 : AO22X1 port map( IN1 => RAM_11_55_port, IN2 => n4533, IN3 => 
                           RAM_10_55_port, IN4 => n4522, Q => n3913);
   U5183 : AO221X1 port map( IN1 => RAM_8_55_port, IN2 => n4555, IN3 => 
                           RAM_9_55_port, IN4 => n4544, IN5 => n3913, Q => 
                           n3920);
   U5184 : AO22X1 port map( IN1 => RAM_15_55_port, IN2 => n4577, IN3 => 
                           RAM_14_55_port, IN4 => n4566, Q => n3914);
   U5185 : AO221X1 port map( IN1 => RAM_12_55_port, IN2 => n4599, IN3 => 
                           RAM_13_55_port, IN4 => n4588, IN5 => n3914, Q => 
                           n3919);
   U5186 : AO22X1 port map( IN1 => RAM_3_55_port, IN2 => n4621, IN3 => 
                           RAM_2_55_port, IN4 => n4610, Q => n3915);
   U5187 : AO221X1 port map( IN1 => RAM_0_55_port, IN2 => n4643, IN3 => 
                           RAM_1_55_port, IN4 => n4632, IN5 => n3915, Q => 
                           n3918);
   U5188 : AO22X1 port map( IN1 => RAM_7_55_port, IN2 => n4665, IN3 => 
                           RAM_6_55_port, IN4 => n4654, Q => n3916);
   U5189 : AO221X1 port map( IN1 => RAM_4_55_port, IN2 => n4687, IN3 => 
                           RAM_5_55_port, IN4 => n4676, IN5 => n3916, Q => 
                           n3917);
   U5190 : OR4X1 port map( IN1 => n3920, IN2 => n3919, IN3 => n3918, IN4 => 
                           n3917, Q => RAMDOUT2(55));
   U5191 : AO22X1 port map( IN1 => RAM_11_56_port, IN2 => n4533, IN3 => 
                           RAM_10_56_port, IN4 => n4522, Q => n3921);
   U5192 : AO221X1 port map( IN1 => RAM_8_56_port, IN2 => n4555, IN3 => 
                           RAM_9_56_port, IN4 => n4544, IN5 => n3921, Q => 
                           n3928);
   U5193 : AO22X1 port map( IN1 => RAM_15_56_port, IN2 => n4577, IN3 => 
                           RAM_14_56_port, IN4 => n4566, Q => n3922);
   U5194 : AO221X1 port map( IN1 => RAM_12_56_port, IN2 => n4599, IN3 => 
                           RAM_13_56_port, IN4 => n4588, IN5 => n3922, Q => 
                           n3927);
   U5195 : AO22X1 port map( IN1 => RAM_3_56_port, IN2 => n4621, IN3 => 
                           RAM_2_56_port, IN4 => n4610, Q => n3923);
   U5196 : AO221X1 port map( IN1 => RAM_0_56_port, IN2 => n4643, IN3 => 
                           RAM_1_56_port, IN4 => n4632, IN5 => n3923, Q => 
                           n3926);
   U5197 : AO22X1 port map( IN1 => RAM_7_56_port, IN2 => n4665, IN3 => 
                           RAM_6_56_port, IN4 => n4654, Q => n3924);
   U5198 : AO221X1 port map( IN1 => RAM_4_56_port, IN2 => n4687, IN3 => 
                           RAM_5_56_port, IN4 => n4676, IN5 => n3924, Q => 
                           n3925);
   U5199 : OR4X1 port map( IN1 => n3928, IN2 => n3927, IN3 => n3926, IN4 => 
                           n3925, Q => RAMDOUT2(56));
   U5200 : AO22X1 port map( IN1 => RAM_11_57_port, IN2 => n4533, IN3 => 
                           RAM_10_57_port, IN4 => n4522, Q => n3929);
   U5201 : AO221X1 port map( IN1 => RAM_8_57_port, IN2 => n4555, IN3 => 
                           RAM_9_57_port, IN4 => n4544, IN5 => n3929, Q => 
                           n3936);
   U5202 : AO22X1 port map( IN1 => RAM_15_57_port, IN2 => n4577, IN3 => 
                           RAM_14_57_port, IN4 => n4566, Q => n3930);
   U5203 : AO221X1 port map( IN1 => RAM_12_57_port, IN2 => n4599, IN3 => 
                           RAM_13_57_port, IN4 => n4588, IN5 => n3930, Q => 
                           n3935);
   U5204 : AO22X1 port map( IN1 => RAM_3_57_port, IN2 => n4621, IN3 => 
                           RAM_2_57_port, IN4 => n4610, Q => n3931);
   U5205 : AO221X1 port map( IN1 => RAM_0_57_port, IN2 => n4643, IN3 => 
                           RAM_1_57_port, IN4 => n4632, IN5 => n3931, Q => 
                           n3934);
   U5206 : AO22X1 port map( IN1 => RAM_7_57_port, IN2 => n4665, IN3 => 
                           RAM_6_57_port, IN4 => n4654, Q => n3932);
   U5207 : AO221X1 port map( IN1 => RAM_4_57_port, IN2 => n4687, IN3 => 
                           RAM_5_57_port, IN4 => n4676, IN5 => n3932, Q => 
                           n3933);
   U5208 : OR4X1 port map( IN1 => n3936, IN2 => n3935, IN3 => n3934, IN4 => 
                           n3933, Q => RAMDOUT2(57));
   U5209 : AO22X1 port map( IN1 => RAM_11_58_port, IN2 => n4533, IN3 => 
                           RAM_10_58_port, IN4 => n4522, Q => n3937);
   U5210 : AO221X1 port map( IN1 => RAM_8_58_port, IN2 => n4555, IN3 => 
                           RAM_9_58_port, IN4 => n4544, IN5 => n3937, Q => 
                           n3944);
   U5211 : AO22X1 port map( IN1 => RAM_15_58_port, IN2 => n4577, IN3 => 
                           RAM_14_58_port, IN4 => n4566, Q => n3938);
   U5212 : AO221X1 port map( IN1 => RAM_12_58_port, IN2 => n4599, IN3 => 
                           RAM_13_58_port, IN4 => n4588, IN5 => n3938, Q => 
                           n3943);
   U5213 : AO22X1 port map( IN1 => RAM_3_58_port, IN2 => n4621, IN3 => 
                           RAM_2_58_port, IN4 => n4610, Q => n3939);
   U5214 : AO221X1 port map( IN1 => RAM_0_58_port, IN2 => n4643, IN3 => 
                           RAM_1_58_port, IN4 => n4632, IN5 => n3939, Q => 
                           n3942);
   U5215 : AO22X1 port map( IN1 => RAM_7_58_port, IN2 => n4665, IN3 => 
                           RAM_6_58_port, IN4 => n4654, Q => n3940);
   U5216 : AO221X1 port map( IN1 => RAM_4_58_port, IN2 => n4687, IN3 => 
                           RAM_5_58_port, IN4 => n4676, IN5 => n3940, Q => 
                           n3941);
   U5217 : OR4X1 port map( IN1 => n3944, IN2 => n3943, IN3 => n3942, IN4 => 
                           n3941, Q => RAMDOUT2(58));
   U5218 : AO22X1 port map( IN1 => RAM_11_59_port, IN2 => n4533, IN3 => 
                           RAM_10_59_port, IN4 => n4522, Q => n3945);
   U5219 : AO221X1 port map( IN1 => RAM_8_59_port, IN2 => n4555, IN3 => 
                           RAM_9_59_port, IN4 => n4544, IN5 => n3945, Q => 
                           n3952);
   U5220 : AO22X1 port map( IN1 => RAM_15_59_port, IN2 => n4577, IN3 => 
                           RAM_14_59_port, IN4 => n4566, Q => n3946);
   U5221 : AO221X1 port map( IN1 => RAM_12_59_port, IN2 => n4599, IN3 => 
                           RAM_13_59_port, IN4 => n4588, IN5 => n3946, Q => 
                           n3951);
   U5222 : AO22X1 port map( IN1 => RAM_3_59_port, IN2 => n4621, IN3 => 
                           RAM_2_59_port, IN4 => n4610, Q => n3947);
   U5223 : AO221X1 port map( IN1 => RAM_0_59_port, IN2 => n4643, IN3 => 
                           RAM_1_59_port, IN4 => n4632, IN5 => n3947, Q => 
                           n3950);
   U5224 : AO22X1 port map( IN1 => RAM_7_59_port, IN2 => n4665, IN3 => 
                           RAM_6_59_port, IN4 => n4654, Q => n3948);
   U5225 : AO221X1 port map( IN1 => RAM_4_59_port, IN2 => n4687, IN3 => 
                           RAM_5_59_port, IN4 => n4676, IN5 => n3948, Q => 
                           n3949);
   U5226 : OR4X1 port map( IN1 => n3952, IN2 => n3951, IN3 => n3950, IN4 => 
                           n3949, Q => RAMDOUT2(59));
   U5227 : AO22X1 port map( IN1 => RAM_11_60_port, IN2 => n4532, IN3 => 
                           RAM_10_60_port, IN4 => n4521, Q => n3953);
   U5228 : AO221X1 port map( IN1 => RAM_8_60_port, IN2 => n4554, IN3 => 
                           RAM_9_60_port, IN4 => n4543, IN5 => n3953, Q => 
                           n3960);
   U5229 : AO22X1 port map( IN1 => RAM_15_60_port, IN2 => n4576, IN3 => 
                           RAM_14_60_port, IN4 => n4565, Q => n3954);
   U5230 : AO221X1 port map( IN1 => RAM_12_60_port, IN2 => n4598, IN3 => 
                           RAM_13_60_port, IN4 => n4587, IN5 => n3954, Q => 
                           n3959);
   U5231 : AO22X1 port map( IN1 => RAM_3_60_port, IN2 => n4620, IN3 => 
                           RAM_2_60_port, IN4 => n4609, Q => n3955);
   U5232 : AO221X1 port map( IN1 => RAM_0_60_port, IN2 => n4642, IN3 => 
                           RAM_1_60_port, IN4 => n4631, IN5 => n3955, Q => 
                           n3958);
   U5233 : AO22X1 port map( IN1 => RAM_7_60_port, IN2 => n4664, IN3 => 
                           RAM_6_60_port, IN4 => n4653, Q => n3956);
   U5234 : AO221X1 port map( IN1 => RAM_4_60_port, IN2 => n4686, IN3 => 
                           RAM_5_60_port, IN4 => n4675, IN5 => n3956, Q => 
                           n3957);
   U5235 : OR4X1 port map( IN1 => n3960, IN2 => n3959, IN3 => n3958, IN4 => 
                           n3957, Q => RAMDOUT2(60));
   U5236 : AO22X1 port map( IN1 => RAM_11_61_port, IN2 => n4532, IN3 => 
                           RAM_10_61_port, IN4 => n4521, Q => n3961);
   U5237 : AO221X1 port map( IN1 => RAM_8_61_port, IN2 => n4554, IN3 => 
                           RAM_9_61_port, IN4 => n4543, IN5 => n3961, Q => 
                           n3968);
   U5238 : AO22X1 port map( IN1 => RAM_15_61_port, IN2 => n4576, IN3 => 
                           RAM_14_61_port, IN4 => n4565, Q => n3962);
   U5239 : AO221X1 port map( IN1 => RAM_12_61_port, IN2 => n4598, IN3 => 
                           RAM_13_61_port, IN4 => n4587, IN5 => n3962, Q => 
                           n3967);
   U5240 : AO22X1 port map( IN1 => RAM_3_61_port, IN2 => n4620, IN3 => 
                           RAM_2_61_port, IN4 => n4609, Q => n3963);
   U5241 : AO221X1 port map( IN1 => RAM_0_61_port, IN2 => n4642, IN3 => 
                           RAM_1_61_port, IN4 => n4631, IN5 => n3963, Q => 
                           n3966);
   U5242 : AO22X1 port map( IN1 => RAM_7_61_port, IN2 => n4664, IN3 => 
                           RAM_6_61_port, IN4 => n4653, Q => n3964);
   U5243 : AO221X1 port map( IN1 => RAM_4_61_port, IN2 => n4686, IN3 => 
                           RAM_5_61_port, IN4 => n4675, IN5 => n3964, Q => 
                           n3965);
   U5244 : OR4X1 port map( IN1 => n3968, IN2 => n3967, IN3 => n3966, IN4 => 
                           n3965, Q => RAMDOUT2(61));
   U5245 : AO22X1 port map( IN1 => RAM_11_62_port, IN2 => n4532, IN3 => 
                           RAM_10_62_port, IN4 => n4521, Q => n3969);
   U5246 : AO221X1 port map( IN1 => RAM_8_62_port, IN2 => n4554, IN3 => 
                           RAM_9_62_port, IN4 => n4543, IN5 => n3969, Q => 
                           n3976);
   U5247 : AO22X1 port map( IN1 => RAM_15_62_port, IN2 => n4576, IN3 => 
                           RAM_14_62_port, IN4 => n4565, Q => n3970);
   U5248 : AO221X1 port map( IN1 => RAM_12_62_port, IN2 => n4598, IN3 => 
                           RAM_13_62_port, IN4 => n4587, IN5 => n3970, Q => 
                           n3975);
   U5249 : AO22X1 port map( IN1 => RAM_3_62_port, IN2 => n4620, IN3 => 
                           RAM_2_62_port, IN4 => n4609, Q => n3971);
   U5250 : AO221X1 port map( IN1 => RAM_0_62_port, IN2 => n4642, IN3 => 
                           RAM_1_62_port, IN4 => n4631, IN5 => n3971, Q => 
                           n3974);
   U5251 : AO22X1 port map( IN1 => RAM_7_62_port, IN2 => n4664, IN3 => 
                           RAM_6_62_port, IN4 => n4653, Q => n3972);
   U5252 : AO221X1 port map( IN1 => RAM_4_62_port, IN2 => n4686, IN3 => 
                           RAM_5_62_port, IN4 => n4675, IN5 => n3972, Q => 
                           n3973);
   U5253 : OR4X1 port map( IN1 => n3976, IN2 => n3975, IN3 => n3974, IN4 => 
                           n3973, Q => RAMDOUT2(62));
   U5254 : AO22X1 port map( IN1 => RAM_11_63_port, IN2 => n4532, IN3 => 
                           RAM_10_63_port, IN4 => n4521, Q => n3977);
   U5255 : AO221X1 port map( IN1 => RAM_8_63_port, IN2 => n4554, IN3 => 
                           RAM_9_63_port, IN4 => n4543, IN5 => n3977, Q => 
                           n3984);
   U5256 : AO22X1 port map( IN1 => RAM_15_63_port, IN2 => n4576, IN3 => 
                           RAM_14_63_port, IN4 => n4565, Q => n3978);
   U5257 : AO221X1 port map( IN1 => RAM_12_63_port, IN2 => n4598, IN3 => 
                           RAM_13_63_port, IN4 => n4587, IN5 => n3978, Q => 
                           n3983);
   U5258 : AO22X1 port map( IN1 => RAM_3_63_port, IN2 => n4620, IN3 => 
                           RAM_2_63_port, IN4 => n4609, Q => n3979);
   U5259 : AO221X1 port map( IN1 => RAM_0_63_port, IN2 => n4642, IN3 => 
                           RAM_1_63_port, IN4 => n4631, IN5 => n3979, Q => 
                           n3982);
   U5260 : AO22X1 port map( IN1 => RAM_7_63_port, IN2 => n4664, IN3 => 
                           RAM_6_63_port, IN4 => n4653, Q => n3980);
   U5261 : AO221X1 port map( IN1 => RAM_4_63_port, IN2 => n4686, IN3 => 
                           RAM_5_63_port, IN4 => n4675, IN5 => n3980, Q => 
                           n3981);
   U5262 : OR4X1 port map( IN1 => n3984, IN2 => n3983, IN3 => n3982, IN4 => 
                           n3981, Q => RAMDOUT2(63));
   U5263 : AO22X1 port map( IN1 => RAM_11_64_port, IN2 => n4532, IN3 => 
                           RAM_10_64_port, IN4 => n4521, Q => n3985);
   U5264 : AO221X1 port map( IN1 => RAM_8_64_port, IN2 => n4554, IN3 => 
                           RAM_9_64_port, IN4 => n4543, IN5 => n3985, Q => 
                           n3992);
   U5265 : AO22X1 port map( IN1 => RAM_15_64_port, IN2 => n4576, IN3 => 
                           RAM_14_64_port, IN4 => n4565, Q => n3986);
   U5266 : AO221X1 port map( IN1 => RAM_12_64_port, IN2 => n4598, IN3 => 
                           RAM_13_64_port, IN4 => n4587, IN5 => n3986, Q => 
                           n3991);
   U5267 : AO22X1 port map( IN1 => RAM_3_64_port, IN2 => n4620, IN3 => 
                           RAM_2_64_port, IN4 => n4609, Q => n3987);
   U5268 : AO221X1 port map( IN1 => RAM_0_64_port, IN2 => n4642, IN3 => 
                           RAM_1_64_port, IN4 => n4631, IN5 => n3987, Q => 
                           n3990);
   U5269 : AO22X1 port map( IN1 => RAM_7_64_port, IN2 => n4664, IN3 => 
                           RAM_6_64_port, IN4 => n4653, Q => n3988);
   U5270 : AO221X1 port map( IN1 => RAM_4_64_port, IN2 => n4686, IN3 => 
                           RAM_5_64_port, IN4 => n4675, IN5 => n3988, Q => 
                           n3989);
   U5271 : OR4X1 port map( IN1 => n3992, IN2 => n3991, IN3 => n3990, IN4 => 
                           n3989, Q => RAMDOUT2(64));
   U5272 : AO22X1 port map( IN1 => RAM_11_65_port, IN2 => n4532, IN3 => 
                           RAM_10_65_port, IN4 => n4521, Q => n3993);
   U5273 : AO221X1 port map( IN1 => RAM_8_65_port, IN2 => n4554, IN3 => 
                           RAM_9_65_port, IN4 => n4543, IN5 => n3993, Q => 
                           n4000);
   U5274 : AO22X1 port map( IN1 => RAM_15_65_port, IN2 => n4576, IN3 => 
                           RAM_14_65_port, IN4 => n4565, Q => n3994);
   U5275 : AO221X1 port map( IN1 => RAM_12_65_port, IN2 => n4598, IN3 => 
                           RAM_13_65_port, IN4 => n4587, IN5 => n3994, Q => 
                           n3999);
   U5276 : AO22X1 port map( IN1 => RAM_3_65_port, IN2 => n4620, IN3 => 
                           RAM_2_65_port, IN4 => n4609, Q => n3995);
   U5277 : AO221X1 port map( IN1 => RAM_0_65_port, IN2 => n4642, IN3 => 
                           RAM_1_65_port, IN4 => n4631, IN5 => n3995, Q => 
                           n3998);
   U5278 : AO22X1 port map( IN1 => RAM_7_65_port, IN2 => n4664, IN3 => 
                           RAM_6_65_port, IN4 => n4653, Q => n3996);
   U5279 : AO221X1 port map( IN1 => RAM_4_65_port, IN2 => n4686, IN3 => 
                           RAM_5_65_port, IN4 => n4675, IN5 => n3996, Q => 
                           n3997);
   U5280 : OR4X1 port map( IN1 => n4000, IN2 => n3999, IN3 => n3998, IN4 => 
                           n3997, Q => RAMDOUT2(65));
   U5281 : AO22X1 port map( IN1 => RAM_11_66_port, IN2 => n4532, IN3 => 
                           RAM_10_66_port, IN4 => n4521, Q => n4001);
   U5282 : AO221X1 port map( IN1 => RAM_8_66_port, IN2 => n4554, IN3 => 
                           RAM_9_66_port, IN4 => n4543, IN5 => n4001, Q => 
                           n4008);
   U5283 : AO22X1 port map( IN1 => RAM_15_66_port, IN2 => n4576, IN3 => 
                           RAM_14_66_port, IN4 => n4565, Q => n4002);
   U5284 : AO221X1 port map( IN1 => RAM_12_66_port, IN2 => n4598, IN3 => 
                           RAM_13_66_port, IN4 => n4587, IN5 => n4002, Q => 
                           n4007);
   U5285 : AO22X1 port map( IN1 => RAM_3_66_port, IN2 => n4620, IN3 => 
                           RAM_2_66_port, IN4 => n4609, Q => n4003);
   U5286 : AO221X1 port map( IN1 => RAM_0_66_port, IN2 => n4642, IN3 => 
                           RAM_1_66_port, IN4 => n4631, IN5 => n4003, Q => 
                           n4006);
   U5287 : AO22X1 port map( IN1 => RAM_7_66_port, IN2 => n4664, IN3 => 
                           RAM_6_66_port, IN4 => n4653, Q => n4004);
   U5288 : AO221X1 port map( IN1 => RAM_4_66_port, IN2 => n4686, IN3 => 
                           RAM_5_66_port, IN4 => n4675, IN5 => n4004, Q => 
                           n4005);
   U5289 : OR4X1 port map( IN1 => n4008, IN2 => n4007, IN3 => n4006, IN4 => 
                           n4005, Q => RAMDOUT2(66));
   U5290 : AO22X1 port map( IN1 => RAM_11_67_port, IN2 => n4532, IN3 => 
                           RAM_10_67_port, IN4 => n4521, Q => n4009);
   U5291 : AO221X1 port map( IN1 => RAM_8_67_port, IN2 => n4554, IN3 => 
                           RAM_9_67_port, IN4 => n4543, IN5 => n4009, Q => 
                           n4016);
   U5292 : AO22X1 port map( IN1 => RAM_15_67_port, IN2 => n4576, IN3 => 
                           RAM_14_67_port, IN4 => n4565, Q => n4010);
   U5293 : AO221X1 port map( IN1 => RAM_12_67_port, IN2 => n4598, IN3 => 
                           RAM_13_67_port, IN4 => n4587, IN5 => n4010, Q => 
                           n4015);
   U5294 : AO22X1 port map( IN1 => RAM_3_67_port, IN2 => n4620, IN3 => 
                           RAM_2_67_port, IN4 => n4609, Q => n4011);
   U5295 : AO221X1 port map( IN1 => RAM_0_67_port, IN2 => n4642, IN3 => 
                           RAM_1_67_port, IN4 => n4631, IN5 => n4011, Q => 
                           n4014);
   U5296 : AO22X1 port map( IN1 => RAM_7_67_port, IN2 => n4664, IN3 => 
                           RAM_6_67_port, IN4 => n4653, Q => n4012);
   U5297 : AO221X1 port map( IN1 => RAM_4_67_port, IN2 => n4686, IN3 => 
                           RAM_5_67_port, IN4 => n4675, IN5 => n4012, Q => 
                           n4013);
   U5298 : OR4X1 port map( IN1 => n4016, IN2 => n4015, IN3 => n4014, IN4 => 
                           n4013, Q => RAMDOUT2(67));
   U5299 : AO22X1 port map( IN1 => RAM_11_68_port, IN2 => n4532, IN3 => 
                           RAM_10_68_port, IN4 => n4521, Q => n4017);
   U5300 : AO221X1 port map( IN1 => RAM_8_68_port, IN2 => n4554, IN3 => 
                           RAM_9_68_port, IN4 => n4543, IN5 => n4017, Q => 
                           n4024);
   U5301 : AO22X1 port map( IN1 => RAM_15_68_port, IN2 => n4576, IN3 => 
                           RAM_14_68_port, IN4 => n4565, Q => n4018);
   U5302 : AO221X1 port map( IN1 => RAM_12_68_port, IN2 => n4598, IN3 => 
                           RAM_13_68_port, IN4 => n4587, IN5 => n4018, Q => 
                           n4023);
   U5303 : AO22X1 port map( IN1 => RAM_3_68_port, IN2 => n4620, IN3 => 
                           RAM_2_68_port, IN4 => n4609, Q => n4019);
   U5304 : AO221X1 port map( IN1 => RAM_0_68_port, IN2 => n4642, IN3 => 
                           RAM_1_68_port, IN4 => n4631, IN5 => n4019, Q => 
                           n4022);
   U5305 : AO22X1 port map( IN1 => RAM_7_68_port, IN2 => n4664, IN3 => 
                           RAM_6_68_port, IN4 => n4653, Q => n4020);
   U5306 : AO221X1 port map( IN1 => RAM_4_68_port, IN2 => n4686, IN3 => 
                           RAM_5_68_port, IN4 => n4675, IN5 => n4020, Q => 
                           n4021);
   U5307 : OR4X1 port map( IN1 => n4024, IN2 => n4023, IN3 => n4022, IN4 => 
                           n4021, Q => RAMDOUT2(68));
   U5308 : AO22X1 port map( IN1 => RAM_11_69_port, IN2 => n4532, IN3 => 
                           RAM_10_69_port, IN4 => n4521, Q => n4025);
   U5309 : AO221X1 port map( IN1 => RAM_8_69_port, IN2 => n4554, IN3 => 
                           RAM_9_69_port, IN4 => n4543, IN5 => n4025, Q => 
                           n4032);
   U5310 : AO22X1 port map( IN1 => RAM_15_69_port, IN2 => n4576, IN3 => 
                           RAM_14_69_port, IN4 => n4565, Q => n4026);
   U5311 : AO221X1 port map( IN1 => RAM_12_69_port, IN2 => n4598, IN3 => 
                           RAM_13_69_port, IN4 => n4587, IN5 => n4026, Q => 
                           n4031);
   U5312 : AO22X1 port map( IN1 => RAM_3_69_port, IN2 => n4620, IN3 => 
                           RAM_2_69_port, IN4 => n4609, Q => n4027);
   U5313 : AO221X1 port map( IN1 => RAM_0_69_port, IN2 => n4642, IN3 => 
                           RAM_1_69_port, IN4 => n4631, IN5 => n4027, Q => 
                           n4030);
   U5314 : AO22X1 port map( IN1 => RAM_7_69_port, IN2 => n4664, IN3 => 
                           RAM_6_69_port, IN4 => n4653, Q => n4028);
   U5315 : AO221X1 port map( IN1 => RAM_4_69_port, IN2 => n4686, IN3 => 
                           RAM_5_69_port, IN4 => n4675, IN5 => n4028, Q => 
                           n4029);
   U5316 : OR4X1 port map( IN1 => n4032, IN2 => n4031, IN3 => n4030, IN4 => 
                           n4029, Q => RAMDOUT2(69));
   U5317 : AO22X1 port map( IN1 => RAM_11_70_port, IN2 => n4532, IN3 => 
                           RAM_10_70_port, IN4 => n4521, Q => n4033);
   U5318 : AO221X1 port map( IN1 => RAM_8_70_port, IN2 => n4554, IN3 => 
                           RAM_9_70_port, IN4 => n4543, IN5 => n4033, Q => 
                           n4040);
   U5319 : AO22X1 port map( IN1 => RAM_15_70_port, IN2 => n4576, IN3 => 
                           RAM_14_70_port, IN4 => n4565, Q => n4034);
   U5320 : AO221X1 port map( IN1 => RAM_12_70_port, IN2 => n4598, IN3 => 
                           RAM_13_70_port, IN4 => n4587, IN5 => n4034, Q => 
                           n4039);
   U5321 : AO22X1 port map( IN1 => RAM_3_70_port, IN2 => n4620, IN3 => 
                           RAM_2_70_port, IN4 => n4609, Q => n4035);
   U5322 : AO221X1 port map( IN1 => RAM_0_70_port, IN2 => n4642, IN3 => 
                           RAM_1_70_port, IN4 => n4631, IN5 => n4035, Q => 
                           n4038);
   U5323 : AO22X1 port map( IN1 => RAM_7_70_port, IN2 => n4664, IN3 => 
                           RAM_6_70_port, IN4 => n4653, Q => n4036);
   U5324 : AO221X1 port map( IN1 => RAM_4_70_port, IN2 => n4686, IN3 => 
                           RAM_5_70_port, IN4 => n4675, IN5 => n4036, Q => 
                           n4037);
   U5325 : OR4X1 port map( IN1 => n4040, IN2 => n4039, IN3 => n4038, IN4 => 
                           n4037, Q => RAMDOUT2(70));
   U5326 : AO22X1 port map( IN1 => RAM_11_71_port, IN2 => n4532, IN3 => 
                           RAM_10_71_port, IN4 => n4521, Q => n4041);
   U5327 : AO221X1 port map( IN1 => RAM_8_71_port, IN2 => n4554, IN3 => 
                           RAM_9_71_port, IN4 => n4543, IN5 => n4041, Q => 
                           n4048);
   U5328 : AO22X1 port map( IN1 => RAM_15_71_port, IN2 => n4576, IN3 => 
                           RAM_14_71_port, IN4 => n4565, Q => n4042);
   U5329 : AO221X1 port map( IN1 => RAM_12_71_port, IN2 => n4598, IN3 => 
                           RAM_13_71_port, IN4 => n4587, IN5 => n4042, Q => 
                           n4047);
   U5330 : AO22X1 port map( IN1 => RAM_3_71_port, IN2 => n4620, IN3 => 
                           RAM_2_71_port, IN4 => n4609, Q => n4043);
   U5331 : AO221X1 port map( IN1 => RAM_0_71_port, IN2 => n4642, IN3 => 
                           RAM_1_71_port, IN4 => n4631, IN5 => n4043, Q => 
                           n4046);
   U5332 : AO22X1 port map( IN1 => RAM_7_71_port, IN2 => n4664, IN3 => 
                           RAM_6_71_port, IN4 => n4653, Q => n4044);
   U5333 : AO221X1 port map( IN1 => RAM_4_71_port, IN2 => n4686, IN3 => 
                           RAM_5_71_port, IN4 => n4675, IN5 => n4044, Q => 
                           n4045);
   U5334 : OR4X1 port map( IN1 => n4048, IN2 => n4047, IN3 => n4046, IN4 => 
                           n4045, Q => RAMDOUT2(71));
   U5335 : AO22X1 port map( IN1 => RAM_11_72_port, IN2 => n4531, IN3 => 
                           RAM_10_72_port, IN4 => n4520, Q => n4049);
   U5336 : AO221X1 port map( IN1 => RAM_8_72_port, IN2 => n4553, IN3 => 
                           RAM_9_72_port, IN4 => n4542, IN5 => n4049, Q => 
                           n4056);
   U5337 : AO22X1 port map( IN1 => RAM_15_72_port, IN2 => n4575, IN3 => 
                           RAM_14_72_port, IN4 => n4564, Q => n4050);
   U5338 : AO221X1 port map( IN1 => RAM_12_72_port, IN2 => n4597, IN3 => 
                           RAM_13_72_port, IN4 => n4586, IN5 => n4050, Q => 
                           n4055);
   U5339 : AO22X1 port map( IN1 => RAM_3_72_port, IN2 => n4619, IN3 => 
                           RAM_2_72_port, IN4 => n4608, Q => n4051);
   U5340 : AO221X1 port map( IN1 => RAM_0_72_port, IN2 => n4641, IN3 => 
                           RAM_1_72_port, IN4 => n4630, IN5 => n4051, Q => 
                           n4054);
   U5341 : AO22X1 port map( IN1 => RAM_7_72_port, IN2 => n4663, IN3 => 
                           RAM_6_72_port, IN4 => n4652, Q => n4052);
   U5342 : AO221X1 port map( IN1 => RAM_4_72_port, IN2 => n4685, IN3 => 
                           RAM_5_72_port, IN4 => n4674, IN5 => n4052, Q => 
                           n4053);
   U5343 : OR4X1 port map( IN1 => n4056, IN2 => n4055, IN3 => n4054, IN4 => 
                           n4053, Q => RAMDOUT2(72));
   U5344 : AO22X1 port map( IN1 => RAM_11_73_port, IN2 => n4531, IN3 => 
                           RAM_10_73_port, IN4 => n4520, Q => n4057);
   U5345 : AO221X1 port map( IN1 => RAM_8_73_port, IN2 => n4553, IN3 => 
                           RAM_9_73_port, IN4 => n4542, IN5 => n4057, Q => 
                           n4064);
   U5346 : AO22X1 port map( IN1 => RAM_15_73_port, IN2 => n4575, IN3 => 
                           RAM_14_73_port, IN4 => n4564, Q => n4058);
   U5347 : AO221X1 port map( IN1 => RAM_12_73_port, IN2 => n4597, IN3 => 
                           RAM_13_73_port, IN4 => n4586, IN5 => n4058, Q => 
                           n4063);
   U5348 : AO22X1 port map( IN1 => RAM_3_73_port, IN2 => n4619, IN3 => 
                           RAM_2_73_port, IN4 => n4608, Q => n4059);
   U5349 : AO221X1 port map( IN1 => RAM_0_73_port, IN2 => n4641, IN3 => 
                           RAM_1_73_port, IN4 => n4630, IN5 => n4059, Q => 
                           n4062);
   U5350 : AO22X1 port map( IN1 => RAM_7_73_port, IN2 => n4663, IN3 => 
                           RAM_6_73_port, IN4 => n4652, Q => n4060);
   U5351 : AO221X1 port map( IN1 => RAM_4_73_port, IN2 => n4685, IN3 => 
                           RAM_5_73_port, IN4 => n4674, IN5 => n4060, Q => 
                           n4061);
   U5352 : OR4X1 port map( IN1 => n4064, IN2 => n4063, IN3 => n4062, IN4 => 
                           n4061, Q => RAMDOUT2(73));
   U5353 : AO22X1 port map( IN1 => RAM_11_74_port, IN2 => n4531, IN3 => 
                           RAM_10_74_port, IN4 => n4520, Q => n4065);
   U5354 : AO221X1 port map( IN1 => RAM_8_74_port, IN2 => n4553, IN3 => 
                           RAM_9_74_port, IN4 => n4542, IN5 => n4065, Q => 
                           n4072);
   U5355 : AO22X1 port map( IN1 => RAM_15_74_port, IN2 => n4575, IN3 => 
                           RAM_14_74_port, IN4 => n4564, Q => n4066);
   U5356 : AO221X1 port map( IN1 => RAM_12_74_port, IN2 => n4597, IN3 => 
                           RAM_13_74_port, IN4 => n4586, IN5 => n4066, Q => 
                           n4071);
   U5357 : AO22X1 port map( IN1 => RAM_3_74_port, IN2 => n4619, IN3 => 
                           RAM_2_74_port, IN4 => n4608, Q => n4067);
   U5358 : AO221X1 port map( IN1 => RAM_0_74_port, IN2 => n4641, IN3 => 
                           RAM_1_74_port, IN4 => n4630, IN5 => n4067, Q => 
                           n4070);
   U5359 : AO22X1 port map( IN1 => RAM_7_74_port, IN2 => n4663, IN3 => 
                           RAM_6_74_port, IN4 => n4652, Q => n4068);
   U5360 : AO221X1 port map( IN1 => RAM_4_74_port, IN2 => n4685, IN3 => 
                           RAM_5_74_port, IN4 => n4674, IN5 => n4068, Q => 
                           n4069);
   U5361 : OR4X1 port map( IN1 => n4072, IN2 => n4071, IN3 => n4070, IN4 => 
                           n4069, Q => RAMDOUT2(74));
   U5362 : AO22X1 port map( IN1 => RAM_11_75_port, IN2 => n4531, IN3 => 
                           RAM_10_75_port, IN4 => n4520, Q => n4073);
   U5363 : AO221X1 port map( IN1 => RAM_8_75_port, IN2 => n4553, IN3 => 
                           RAM_9_75_port, IN4 => n4542, IN5 => n4073, Q => 
                           n4080);
   U5364 : AO22X1 port map( IN1 => RAM_15_75_port, IN2 => n4575, IN3 => 
                           RAM_14_75_port, IN4 => n4564, Q => n4074);
   U5365 : AO221X1 port map( IN1 => RAM_12_75_port, IN2 => n4597, IN3 => 
                           RAM_13_75_port, IN4 => n4586, IN5 => n4074, Q => 
                           n4079);
   U5366 : AO22X1 port map( IN1 => RAM_3_75_port, IN2 => n4619, IN3 => 
                           RAM_2_75_port, IN4 => n4608, Q => n4075);
   U5367 : AO221X1 port map( IN1 => RAM_0_75_port, IN2 => n4641, IN3 => 
                           RAM_1_75_port, IN4 => n4630, IN5 => n4075, Q => 
                           n4078);
   U5368 : AO22X1 port map( IN1 => RAM_7_75_port, IN2 => n4663, IN3 => 
                           RAM_6_75_port, IN4 => n4652, Q => n4076);
   U5369 : AO221X1 port map( IN1 => RAM_4_75_port, IN2 => n4685, IN3 => 
                           RAM_5_75_port, IN4 => n4674, IN5 => n4076, Q => 
                           n4077);
   U5370 : OR4X1 port map( IN1 => n4080, IN2 => n4079, IN3 => n4078, IN4 => 
                           n4077, Q => RAMDOUT2(75));
   U5371 : AO22X1 port map( IN1 => RAM_11_76_port, IN2 => n4531, IN3 => 
                           RAM_10_76_port, IN4 => n4520, Q => n4081);
   U5372 : AO221X1 port map( IN1 => RAM_8_76_port, IN2 => n4553, IN3 => 
                           RAM_9_76_port, IN4 => n4542, IN5 => n4081, Q => 
                           n4088);
   U5373 : AO22X1 port map( IN1 => RAM_15_76_port, IN2 => n4575, IN3 => 
                           RAM_14_76_port, IN4 => n4564, Q => n4082);
   U5374 : AO221X1 port map( IN1 => RAM_12_76_port, IN2 => n4597, IN3 => 
                           RAM_13_76_port, IN4 => n4586, IN5 => n4082, Q => 
                           n4087);
   U5375 : AO22X1 port map( IN1 => RAM_3_76_port, IN2 => n4619, IN3 => 
                           RAM_2_76_port, IN4 => n4608, Q => n4083);
   U5376 : AO221X1 port map( IN1 => RAM_0_76_port, IN2 => n4641, IN3 => 
                           RAM_1_76_port, IN4 => n4630, IN5 => n4083, Q => 
                           n4086);
   U5377 : AO22X1 port map( IN1 => RAM_7_76_port, IN2 => n4663, IN3 => 
                           RAM_6_76_port, IN4 => n4652, Q => n4084);
   U5378 : AO221X1 port map( IN1 => RAM_4_76_port, IN2 => n4685, IN3 => 
                           RAM_5_76_port, IN4 => n4674, IN5 => n4084, Q => 
                           n4085);
   U5379 : OR4X1 port map( IN1 => n4088, IN2 => n4087, IN3 => n4086, IN4 => 
                           n4085, Q => RAMDOUT2(76));
   U5380 : AO22X1 port map( IN1 => RAM_11_77_port, IN2 => n4531, IN3 => 
                           RAM_10_77_port, IN4 => n4520, Q => n4089);
   U5381 : AO221X1 port map( IN1 => RAM_8_77_port, IN2 => n4553, IN3 => 
                           RAM_9_77_port, IN4 => n4542, IN5 => n4089, Q => 
                           n4096);
   U5382 : AO22X1 port map( IN1 => RAM_15_77_port, IN2 => n4575, IN3 => 
                           RAM_14_77_port, IN4 => n4564, Q => n4090);
   U5383 : AO221X1 port map( IN1 => RAM_12_77_port, IN2 => n4597, IN3 => 
                           RAM_13_77_port, IN4 => n4586, IN5 => n4090, Q => 
                           n4095);
   U5384 : AO22X1 port map( IN1 => RAM_3_77_port, IN2 => n4619, IN3 => 
                           RAM_2_77_port, IN4 => n4608, Q => n4091);
   U5385 : AO221X1 port map( IN1 => RAM_0_77_port, IN2 => n4641, IN3 => 
                           RAM_1_77_port, IN4 => n4630, IN5 => n4091, Q => 
                           n4094);
   U5386 : AO22X1 port map( IN1 => RAM_7_77_port, IN2 => n4663, IN3 => 
                           RAM_6_77_port, IN4 => n4652, Q => n4092);
   U5387 : AO221X1 port map( IN1 => RAM_4_77_port, IN2 => n4685, IN3 => 
                           RAM_5_77_port, IN4 => n4674, IN5 => n4092, Q => 
                           n4093);
   U5388 : OR4X1 port map( IN1 => n4096, IN2 => n4095, IN3 => n4094, IN4 => 
                           n4093, Q => RAMDOUT2(77));
   U5389 : AO22X1 port map( IN1 => RAM_11_78_port, IN2 => n4531, IN3 => 
                           RAM_10_78_port, IN4 => n4520, Q => n4097);
   U5390 : AO221X1 port map( IN1 => RAM_8_78_port, IN2 => n4553, IN3 => 
                           RAM_9_78_port, IN4 => n4542, IN5 => n4097, Q => 
                           n4104);
   U5391 : AO22X1 port map( IN1 => RAM_15_78_port, IN2 => n4575, IN3 => 
                           RAM_14_78_port, IN4 => n4564, Q => n4098);
   U5392 : AO221X1 port map( IN1 => RAM_12_78_port, IN2 => n4597, IN3 => 
                           RAM_13_78_port, IN4 => n4586, IN5 => n4098, Q => 
                           n4103);
   U5393 : AO22X1 port map( IN1 => RAM_3_78_port, IN2 => n4619, IN3 => 
                           RAM_2_78_port, IN4 => n4608, Q => n4099);
   U5394 : AO221X1 port map( IN1 => RAM_0_78_port, IN2 => n4641, IN3 => 
                           RAM_1_78_port, IN4 => n4630, IN5 => n4099, Q => 
                           n4102);
   U5395 : AO22X1 port map( IN1 => RAM_7_78_port, IN2 => n4663, IN3 => 
                           RAM_6_78_port, IN4 => n4652, Q => n4100);
   U5396 : AO221X1 port map( IN1 => RAM_4_78_port, IN2 => n4685, IN3 => 
                           RAM_5_78_port, IN4 => n4674, IN5 => n4100, Q => 
                           n4101);
   U5397 : OR4X1 port map( IN1 => n4104, IN2 => n4103, IN3 => n4102, IN4 => 
                           n4101, Q => RAMDOUT2(78));
   U5398 : AO22X1 port map( IN1 => RAM_11_79_port, IN2 => n4531, IN3 => 
                           RAM_10_79_port, IN4 => n4520, Q => n4105);
   U5399 : AO221X1 port map( IN1 => RAM_8_79_port, IN2 => n4553, IN3 => 
                           RAM_9_79_port, IN4 => n4542, IN5 => n4105, Q => 
                           n4112);
   U5400 : AO22X1 port map( IN1 => RAM_15_79_port, IN2 => n4575, IN3 => 
                           RAM_14_79_port, IN4 => n4564, Q => n4106);
   U5401 : AO221X1 port map( IN1 => RAM_12_79_port, IN2 => n4597, IN3 => 
                           RAM_13_79_port, IN4 => n4586, IN5 => n4106, Q => 
                           n4111);
   U5402 : AO22X1 port map( IN1 => RAM_3_79_port, IN2 => n4619, IN3 => 
                           RAM_2_79_port, IN4 => n4608, Q => n4107);
   U5403 : AO221X1 port map( IN1 => RAM_0_79_port, IN2 => n4641, IN3 => 
                           RAM_1_79_port, IN4 => n4630, IN5 => n4107, Q => 
                           n4110);
   U5404 : AO22X1 port map( IN1 => RAM_7_79_port, IN2 => n4663, IN3 => 
                           RAM_6_79_port, IN4 => n4652, Q => n4108);
   U5405 : AO221X1 port map( IN1 => RAM_4_79_port, IN2 => n4685, IN3 => 
                           RAM_5_79_port, IN4 => n4674, IN5 => n4108, Q => 
                           n4109);
   U5406 : OR4X1 port map( IN1 => n4112, IN2 => n4111, IN3 => n4110, IN4 => 
                           n4109, Q => RAMDOUT2(79));
   U5407 : AO22X1 port map( IN1 => RAM_11_80_port, IN2 => n4531, IN3 => 
                           RAM_10_80_port, IN4 => n4520, Q => n4113);
   U5408 : AO221X1 port map( IN1 => RAM_8_80_port, IN2 => n4553, IN3 => 
                           RAM_9_80_port, IN4 => n4542, IN5 => n4113, Q => 
                           n4120);
   U5409 : AO22X1 port map( IN1 => RAM_15_80_port, IN2 => n4575, IN3 => 
                           RAM_14_80_port, IN4 => n4564, Q => n4114);
   U5410 : AO221X1 port map( IN1 => RAM_12_80_port, IN2 => n4597, IN3 => 
                           RAM_13_80_port, IN4 => n4586, IN5 => n4114, Q => 
                           n4119);
   U5411 : AO22X1 port map( IN1 => RAM_3_80_port, IN2 => n4619, IN3 => 
                           RAM_2_80_port, IN4 => n4608, Q => n4115);
   U5412 : AO221X1 port map( IN1 => RAM_0_80_port, IN2 => n4641, IN3 => 
                           RAM_1_80_port, IN4 => n4630, IN5 => n4115, Q => 
                           n4118);
   U5413 : AO22X1 port map( IN1 => RAM_7_80_port, IN2 => n4663, IN3 => 
                           RAM_6_80_port, IN4 => n4652, Q => n4116);
   U5414 : AO221X1 port map( IN1 => RAM_4_80_port, IN2 => n4685, IN3 => 
                           RAM_5_80_port, IN4 => n4674, IN5 => n4116, Q => 
                           n4117);
   U5415 : OR4X1 port map( IN1 => n4120, IN2 => n4119, IN3 => n4118, IN4 => 
                           n4117, Q => RAMDOUT2(80));
   U5416 : AO22X1 port map( IN1 => RAM_11_81_port, IN2 => n4531, IN3 => 
                           RAM_10_81_port, IN4 => n4520, Q => n4121);
   U5417 : AO221X1 port map( IN1 => RAM_8_81_port, IN2 => n4553, IN3 => 
                           RAM_9_81_port, IN4 => n4542, IN5 => n4121, Q => 
                           n4128);
   U5418 : AO22X1 port map( IN1 => RAM_15_81_port, IN2 => n4575, IN3 => 
                           RAM_14_81_port, IN4 => n4564, Q => n4122);
   U5419 : AO221X1 port map( IN1 => RAM_12_81_port, IN2 => n4597, IN3 => 
                           RAM_13_81_port, IN4 => n4586, IN5 => n4122, Q => 
                           n4127);
   U5420 : AO22X1 port map( IN1 => RAM_3_81_port, IN2 => n4619, IN3 => 
                           RAM_2_81_port, IN4 => n4608, Q => n4123);
   U5421 : AO221X1 port map( IN1 => RAM_0_81_port, IN2 => n4641, IN3 => 
                           RAM_1_81_port, IN4 => n4630, IN5 => n4123, Q => 
                           n4126);
   U5422 : AO22X1 port map( IN1 => RAM_7_81_port, IN2 => n4663, IN3 => 
                           RAM_6_81_port, IN4 => n4652, Q => n4124);
   U5423 : AO221X1 port map( IN1 => RAM_4_81_port, IN2 => n4685, IN3 => 
                           RAM_5_81_port, IN4 => n4674, IN5 => n4124, Q => 
                           n4125);
   U5424 : OR4X1 port map( IN1 => n4128, IN2 => n4127, IN3 => n4126, IN4 => 
                           n4125, Q => RAMDOUT2(81));
   U5425 : AO22X1 port map( IN1 => RAM_11_82_port, IN2 => n4531, IN3 => 
                           RAM_10_82_port, IN4 => n4520, Q => n4129);
   U5426 : AO221X1 port map( IN1 => RAM_8_82_port, IN2 => n4553, IN3 => 
                           RAM_9_82_port, IN4 => n4542, IN5 => n4129, Q => 
                           n4136);
   U5427 : AO22X1 port map( IN1 => RAM_15_82_port, IN2 => n4575, IN3 => 
                           RAM_14_82_port, IN4 => n4564, Q => n4130);
   U5428 : AO221X1 port map( IN1 => RAM_12_82_port, IN2 => n4597, IN3 => 
                           RAM_13_82_port, IN4 => n4586, IN5 => n4130, Q => 
                           n4135);
   U5429 : AO22X1 port map( IN1 => RAM_3_82_port, IN2 => n4619, IN3 => 
                           RAM_2_82_port, IN4 => n4608, Q => n4131);
   U5430 : AO221X1 port map( IN1 => RAM_0_82_port, IN2 => n4641, IN3 => 
                           RAM_1_82_port, IN4 => n4630, IN5 => n4131, Q => 
                           n4134);
   U5431 : AO22X1 port map( IN1 => RAM_7_82_port, IN2 => n4663, IN3 => 
                           RAM_6_82_port, IN4 => n4652, Q => n4132);
   U5432 : AO221X1 port map( IN1 => RAM_4_82_port, IN2 => n4685, IN3 => 
                           RAM_5_82_port, IN4 => n4674, IN5 => n4132, Q => 
                           n4133);
   U5433 : OR4X1 port map( IN1 => n4136, IN2 => n4135, IN3 => n4134, IN4 => 
                           n4133, Q => RAMDOUT2(82));
   U5434 : AO22X1 port map( IN1 => RAM_11_83_port, IN2 => n4531, IN3 => 
                           RAM_10_83_port, IN4 => n4520, Q => n4137);
   U5435 : AO221X1 port map( IN1 => RAM_8_83_port, IN2 => n4553, IN3 => 
                           RAM_9_83_port, IN4 => n4542, IN5 => n4137, Q => 
                           n4144);
   U5436 : AO22X1 port map( IN1 => RAM_15_83_port, IN2 => n4575, IN3 => 
                           RAM_14_83_port, IN4 => n4564, Q => n4138);
   U5437 : AO221X1 port map( IN1 => RAM_12_83_port, IN2 => n4597, IN3 => 
                           RAM_13_83_port, IN4 => n4586, IN5 => n4138, Q => 
                           n4143);
   U5438 : AO22X1 port map( IN1 => RAM_3_83_port, IN2 => n4619, IN3 => 
                           RAM_2_83_port, IN4 => n4608, Q => n4139);
   U5439 : AO221X1 port map( IN1 => RAM_0_83_port, IN2 => n4641, IN3 => 
                           RAM_1_83_port, IN4 => n4630, IN5 => n4139, Q => 
                           n4142);
   U5440 : AO22X1 port map( IN1 => RAM_7_83_port, IN2 => n4663, IN3 => 
                           RAM_6_83_port, IN4 => n4652, Q => n4140);
   U5441 : AO221X1 port map( IN1 => RAM_4_83_port, IN2 => n4685, IN3 => 
                           RAM_5_83_port, IN4 => n4674, IN5 => n4140, Q => 
                           n4141);
   U5442 : OR4X1 port map( IN1 => n4144, IN2 => n4143, IN3 => n4142, IN4 => 
                           n4141, Q => RAMDOUT2(83));
   U5443 : AO22X1 port map( IN1 => RAM_11_84_port, IN2 => n4530, IN3 => 
                           RAM_10_84_port, IN4 => n4519, Q => n4145);
   U5444 : AO221X1 port map( IN1 => RAM_8_84_port, IN2 => n4552, IN3 => 
                           RAM_9_84_port, IN4 => n4541, IN5 => n4145, Q => 
                           n4152);
   U5445 : AO22X1 port map( IN1 => RAM_15_84_port, IN2 => n4574, IN3 => 
                           RAM_14_84_port, IN4 => n4563, Q => n4146);
   U5446 : AO221X1 port map( IN1 => RAM_12_84_port, IN2 => n4596, IN3 => 
                           RAM_13_84_port, IN4 => n4585, IN5 => n4146, Q => 
                           n4151);
   U5447 : AO22X1 port map( IN1 => RAM_3_84_port, IN2 => n4618, IN3 => 
                           RAM_2_84_port, IN4 => n4607, Q => n4147);
   U5448 : AO221X1 port map( IN1 => RAM_0_84_port, IN2 => n4640, IN3 => 
                           RAM_1_84_port, IN4 => n4629, IN5 => n4147, Q => 
                           n4150);
   U5449 : AO22X1 port map( IN1 => RAM_7_84_port, IN2 => n4662, IN3 => 
                           RAM_6_84_port, IN4 => n4651, Q => n4148);
   U5450 : AO221X1 port map( IN1 => RAM_4_84_port, IN2 => n4684, IN3 => 
                           RAM_5_84_port, IN4 => n4673, IN5 => n4148, Q => 
                           n4149);
   U5451 : OR4X1 port map( IN1 => n4152, IN2 => n4151, IN3 => n4150, IN4 => 
                           n4149, Q => RAMDOUT2(84));
   U5452 : AO22X1 port map( IN1 => RAM_11_85_port, IN2 => n4530, IN3 => 
                           RAM_10_85_port, IN4 => n4519, Q => n4153);
   U5453 : AO221X1 port map( IN1 => RAM_8_85_port, IN2 => n4552, IN3 => 
                           RAM_9_85_port, IN4 => n4541, IN5 => n4153, Q => 
                           n4160);
   U5454 : AO22X1 port map( IN1 => RAM_15_85_port, IN2 => n4574, IN3 => 
                           RAM_14_85_port, IN4 => n4563, Q => n4154);
   U5455 : AO221X1 port map( IN1 => RAM_12_85_port, IN2 => n4596, IN3 => 
                           RAM_13_85_port, IN4 => n4585, IN5 => n4154, Q => 
                           n4159);
   U5456 : AO22X1 port map( IN1 => RAM_3_85_port, IN2 => n4618, IN3 => 
                           RAM_2_85_port, IN4 => n4607, Q => n4155);
   U5457 : AO221X1 port map( IN1 => RAM_0_85_port, IN2 => n4640, IN3 => 
                           RAM_1_85_port, IN4 => n4629, IN5 => n4155, Q => 
                           n4158);
   U5458 : AO22X1 port map( IN1 => RAM_7_85_port, IN2 => n4662, IN3 => 
                           RAM_6_85_port, IN4 => n4651, Q => n4156);
   U5459 : AO221X1 port map( IN1 => RAM_4_85_port, IN2 => n4684, IN3 => 
                           RAM_5_85_port, IN4 => n4673, IN5 => n4156, Q => 
                           n4157);
   U5460 : OR4X1 port map( IN1 => n4160, IN2 => n4159, IN3 => n4158, IN4 => 
                           n4157, Q => RAMDOUT2(85));
   U5461 : AO22X1 port map( IN1 => RAM_11_86_port, IN2 => n4530, IN3 => 
                           RAM_10_86_port, IN4 => n4519, Q => n4161);
   U5462 : AO221X1 port map( IN1 => RAM_8_86_port, IN2 => n4552, IN3 => 
                           RAM_9_86_port, IN4 => n4541, IN5 => n4161, Q => 
                           n4168);
   U5463 : AO22X1 port map( IN1 => RAM_15_86_port, IN2 => n4574, IN3 => 
                           RAM_14_86_port, IN4 => n4563, Q => n4162);
   U5464 : AO221X1 port map( IN1 => RAM_12_86_port, IN2 => n4596, IN3 => 
                           RAM_13_86_port, IN4 => n4585, IN5 => n4162, Q => 
                           n4167);
   U5465 : AO22X1 port map( IN1 => RAM_3_86_port, IN2 => n4618, IN3 => 
                           RAM_2_86_port, IN4 => n4607, Q => n4163);
   U5466 : AO221X1 port map( IN1 => RAM_0_86_port, IN2 => n4640, IN3 => 
                           RAM_1_86_port, IN4 => n4629, IN5 => n4163, Q => 
                           n4166);
   U5467 : AO22X1 port map( IN1 => RAM_7_86_port, IN2 => n4662, IN3 => 
                           RAM_6_86_port, IN4 => n4651, Q => n4164);
   U5468 : AO221X1 port map( IN1 => RAM_4_86_port, IN2 => n4684, IN3 => 
                           RAM_5_86_port, IN4 => n4673, IN5 => n4164, Q => 
                           n4165);
   U5469 : OR4X1 port map( IN1 => n4168, IN2 => n4167, IN3 => n4166, IN4 => 
                           n4165, Q => RAMDOUT2(86));
   U5470 : AO22X1 port map( IN1 => RAM_11_87_port, IN2 => n4530, IN3 => 
                           RAM_10_87_port, IN4 => n4519, Q => n4169);
   U5471 : AO221X1 port map( IN1 => RAM_8_87_port, IN2 => n4552, IN3 => 
                           RAM_9_87_port, IN4 => n4541, IN5 => n4169, Q => 
                           n4176);
   U5472 : AO22X1 port map( IN1 => RAM_15_87_port, IN2 => n4574, IN3 => 
                           RAM_14_87_port, IN4 => n4563, Q => n4170);
   U5473 : AO221X1 port map( IN1 => RAM_12_87_port, IN2 => n4596, IN3 => 
                           RAM_13_87_port, IN4 => n4585, IN5 => n4170, Q => 
                           n4175);
   U5474 : AO22X1 port map( IN1 => RAM_3_87_port, IN2 => n4618, IN3 => 
                           RAM_2_87_port, IN4 => n4607, Q => n4171);
   U5475 : AO221X1 port map( IN1 => RAM_0_87_port, IN2 => n4640, IN3 => 
                           RAM_1_87_port, IN4 => n4629, IN5 => n4171, Q => 
                           n4174);
   U5476 : AO22X1 port map( IN1 => RAM_7_87_port, IN2 => n4662, IN3 => 
                           RAM_6_87_port, IN4 => n4651, Q => n4172);
   U5477 : AO221X1 port map( IN1 => RAM_4_87_port, IN2 => n4684, IN3 => 
                           RAM_5_87_port, IN4 => n4673, IN5 => n4172, Q => 
                           n4173);
   U5478 : OR4X1 port map( IN1 => n4176, IN2 => n4175, IN3 => n4174, IN4 => 
                           n4173, Q => RAMDOUT2(87));
   U5479 : AO22X1 port map( IN1 => RAM_11_88_port, IN2 => n4530, IN3 => 
                           RAM_10_88_port, IN4 => n4519, Q => n4177);
   U5480 : AO221X1 port map( IN1 => RAM_8_88_port, IN2 => n4552, IN3 => 
                           RAM_9_88_port, IN4 => n4541, IN5 => n4177, Q => 
                           n4184);
   U5481 : AO22X1 port map( IN1 => RAM_15_88_port, IN2 => n4574, IN3 => 
                           RAM_14_88_port, IN4 => n4563, Q => n4178);
   U5482 : AO221X1 port map( IN1 => RAM_12_88_port, IN2 => n4596, IN3 => 
                           RAM_13_88_port, IN4 => n4585, IN5 => n4178, Q => 
                           n4183);
   U5483 : AO22X1 port map( IN1 => RAM_3_88_port, IN2 => n4618, IN3 => 
                           RAM_2_88_port, IN4 => n4607, Q => n4179);
   U5484 : AO221X1 port map( IN1 => RAM_0_88_port, IN2 => n4640, IN3 => 
                           RAM_1_88_port, IN4 => n4629, IN5 => n4179, Q => 
                           n4182);
   U5485 : AO22X1 port map( IN1 => RAM_7_88_port, IN2 => n4662, IN3 => 
                           RAM_6_88_port, IN4 => n4651, Q => n4180);
   U5486 : AO221X1 port map( IN1 => RAM_4_88_port, IN2 => n4684, IN3 => 
                           RAM_5_88_port, IN4 => n4673, IN5 => n4180, Q => 
                           n4181);
   U5487 : AO22X1 port map( IN1 => RAM_11_89_port, IN2 => n4530, IN3 => 
                           RAM_10_89_port, IN4 => n4519, Q => n4185);
   U5488 : AO221X1 port map( IN1 => RAM_8_89_port, IN2 => n4552, IN3 => 
                           RAM_9_89_port, IN4 => n4541, IN5 => n4185, Q => 
                           n4192);
   U5489 : AO22X1 port map( IN1 => RAM_15_89_port, IN2 => n4574, IN3 => 
                           RAM_14_89_port, IN4 => n4563, Q => n4186);
   U5490 : AO221X1 port map( IN1 => RAM_12_89_port, IN2 => n4596, IN3 => 
                           RAM_13_89_port, IN4 => n4585, IN5 => n4186, Q => 
                           n4191);
   U5491 : AO22X1 port map( IN1 => RAM_3_89_port, IN2 => n4618, IN3 => 
                           RAM_2_89_port, IN4 => n4607, Q => n4187);
   U5492 : AO221X1 port map( IN1 => RAM_0_89_port, IN2 => n4640, IN3 => 
                           RAM_1_89_port, IN4 => n4629, IN5 => n4187, Q => 
                           n4190);
   U5493 : AO22X1 port map( IN1 => RAM_7_89_port, IN2 => n4662, IN3 => 
                           RAM_6_89_port, IN4 => n4651, Q => n4188);
   U5494 : AO221X1 port map( IN1 => RAM_4_89_port, IN2 => n4684, IN3 => 
                           RAM_5_89_port, IN4 => n4673, IN5 => n4188, Q => 
                           n4189);
   U5495 : OR4X1 port map( IN1 => n4192, IN2 => n4191, IN3 => n4190, IN4 => 
                           n4189, Q => RAMDOUT2(89));
   U5496 : AO22X1 port map( IN1 => RAM_11_90_port, IN2 => n4530, IN3 => 
                           RAM_10_90_port, IN4 => n4519, Q => n4193);
   U5497 : AO221X1 port map( IN1 => RAM_8_90_port, IN2 => n4552, IN3 => 
                           RAM_9_90_port, IN4 => n4541, IN5 => n4193, Q => 
                           n4200);
   U5498 : AO22X1 port map( IN1 => RAM_15_90_port, IN2 => n4574, IN3 => 
                           RAM_14_90_port, IN4 => n4563, Q => n4194);
   U5499 : AO221X1 port map( IN1 => RAM_12_90_port, IN2 => n4596, IN3 => 
                           RAM_13_90_port, IN4 => n4585, IN5 => n4194, Q => 
                           n4199);
   U5500 : AO22X1 port map( IN1 => RAM_3_90_port, IN2 => n4618, IN3 => 
                           RAM_2_90_port, IN4 => n4607, Q => n4195);
   U5501 : AO221X1 port map( IN1 => RAM_0_90_port, IN2 => n4640, IN3 => 
                           RAM_1_90_port, IN4 => n4629, IN5 => n4195, Q => 
                           n4198);
   U5502 : AO22X1 port map( IN1 => RAM_7_90_port, IN2 => n4662, IN3 => 
                           RAM_6_90_port, IN4 => n4651, Q => n4196);
   U5503 : AO221X1 port map( IN1 => RAM_4_90_port, IN2 => n4684, IN3 => 
                           RAM_5_90_port, IN4 => n4673, IN5 => n4196, Q => 
                           n4197);
   U5504 : OR4X1 port map( IN1 => n4200, IN2 => n4199, IN3 => n4198, IN4 => 
                           n4197, Q => RAMDOUT2(90));
   U5505 : AO22X1 port map( IN1 => RAM_11_91_port, IN2 => n4530, IN3 => 
                           RAM_10_91_port, IN4 => n4519, Q => n4201);
   U5506 : AO221X1 port map( IN1 => RAM_8_91_port, IN2 => n4552, IN3 => 
                           RAM_9_91_port, IN4 => n4541, IN5 => n4201, Q => 
                           n4208);
   U5507 : AO22X1 port map( IN1 => RAM_15_91_port, IN2 => n4574, IN3 => 
                           RAM_14_91_port, IN4 => n4563, Q => n4202);
   U5508 : AO221X1 port map( IN1 => RAM_12_91_port, IN2 => n4596, IN3 => 
                           RAM_13_91_port, IN4 => n4585, IN5 => n4202, Q => 
                           n4207);
   U5509 : AO22X1 port map( IN1 => RAM_3_91_port, IN2 => n4618, IN3 => 
                           RAM_2_91_port, IN4 => n4607, Q => n4203);
   U5510 : AO221X1 port map( IN1 => RAM_0_91_port, IN2 => n4640, IN3 => 
                           RAM_1_91_port, IN4 => n4629, IN5 => n4203, Q => 
                           n4206);
   U5511 : AO22X1 port map( IN1 => RAM_7_91_port, IN2 => n4662, IN3 => 
                           RAM_6_91_port, IN4 => n4651, Q => n4204);
   U5512 : AO221X1 port map( IN1 => RAM_4_91_port, IN2 => n4684, IN3 => 
                           RAM_5_91_port, IN4 => n4673, IN5 => n4204, Q => 
                           n4205);
   U5513 : OR4X1 port map( IN1 => n4208, IN2 => n4207, IN3 => n4206, IN4 => 
                           n4205, Q => RAMDOUT2(91));
   U5514 : AO22X1 port map( IN1 => RAM_11_92_port, IN2 => n4530, IN3 => 
                           RAM_10_92_port, IN4 => n4519, Q => n4209);
   U5515 : AO221X1 port map( IN1 => RAM_8_92_port, IN2 => n4552, IN3 => 
                           RAM_9_92_port, IN4 => n4541, IN5 => n4209, Q => 
                           n4216);
   U5516 : AO22X1 port map( IN1 => RAM_15_92_port, IN2 => n4574, IN3 => 
                           RAM_14_92_port, IN4 => n4563, Q => n4210);
   U5517 : AO221X1 port map( IN1 => RAM_12_92_port, IN2 => n4596, IN3 => 
                           RAM_13_92_port, IN4 => n4585, IN5 => n4210, Q => 
                           n4215);
   U5518 : AO22X1 port map( IN1 => RAM_3_92_port, IN2 => n4618, IN3 => 
                           RAM_2_92_port, IN4 => n4607, Q => n4211);
   U5519 : AO221X1 port map( IN1 => RAM_0_92_port, IN2 => n4640, IN3 => 
                           RAM_1_92_port, IN4 => n4629, IN5 => n4211, Q => 
                           n4214);
   U5520 : AO22X1 port map( IN1 => RAM_7_92_port, IN2 => n4662, IN3 => 
                           RAM_6_92_port, IN4 => n4651, Q => n4212);
   U5521 : AO221X1 port map( IN1 => RAM_4_92_port, IN2 => n4684, IN3 => 
                           RAM_5_92_port, IN4 => n4673, IN5 => n4212, Q => 
                           n4213);
   U5522 : OR4X1 port map( IN1 => n4216, IN2 => n4215, IN3 => n4214, IN4 => 
                           n4213, Q => RAMDOUT2(92));
   U5523 : AO22X1 port map( IN1 => RAM_11_93_port, IN2 => n4530, IN3 => 
                           RAM_10_93_port, IN4 => n4519, Q => n4217);
   U5524 : AO221X1 port map( IN1 => RAM_8_93_port, IN2 => n4552, IN3 => 
                           RAM_9_93_port, IN4 => n4541, IN5 => n4217, Q => 
                           n4224);
   U5525 : AO22X1 port map( IN1 => RAM_15_93_port, IN2 => n4574, IN3 => 
                           RAM_14_93_port, IN4 => n4563, Q => n4218);
   U5526 : AO221X1 port map( IN1 => RAM_12_93_port, IN2 => n4596, IN3 => 
                           RAM_13_93_port, IN4 => n4585, IN5 => n4218, Q => 
                           n4223);
   U5527 : AO22X1 port map( IN1 => RAM_3_93_port, IN2 => n4618, IN3 => 
                           RAM_2_93_port, IN4 => n4607, Q => n4219);
   U5528 : AO221X1 port map( IN1 => RAM_0_93_port, IN2 => n4640, IN3 => 
                           RAM_1_93_port, IN4 => n4629, IN5 => n4219, Q => 
                           n4222);
   U5529 : AO22X1 port map( IN1 => RAM_7_93_port, IN2 => n4662, IN3 => 
                           RAM_6_93_port, IN4 => n4651, Q => n4220);
   U5530 : AO221X1 port map( IN1 => RAM_4_93_port, IN2 => n4684, IN3 => 
                           RAM_5_93_port, IN4 => n4673, IN5 => n4220, Q => 
                           n4221);
   U5531 : OR4X1 port map( IN1 => n4224, IN2 => n4223, IN3 => n4222, IN4 => 
                           n4221, Q => RAMDOUT2(93));
   U5532 : AO22X1 port map( IN1 => RAM_11_94_port, IN2 => n4530, IN3 => 
                           RAM_10_94_port, IN4 => n4519, Q => n4225);
   U5533 : AO221X1 port map( IN1 => RAM_8_94_port, IN2 => n4552, IN3 => 
                           RAM_9_94_port, IN4 => n4541, IN5 => n4225, Q => 
                           n4232);
   U5534 : AO22X1 port map( IN1 => RAM_15_94_port, IN2 => n4574, IN3 => 
                           RAM_14_94_port, IN4 => n4563, Q => n4226);
   U5535 : AO221X1 port map( IN1 => RAM_12_94_port, IN2 => n4596, IN3 => 
                           RAM_13_94_port, IN4 => n4585, IN5 => n4226, Q => 
                           n4231);
   U5536 : AO22X1 port map( IN1 => RAM_3_94_port, IN2 => n4618, IN3 => 
                           RAM_2_94_port, IN4 => n4607, Q => n4227);
   U5537 : AO221X1 port map( IN1 => RAM_0_94_port, IN2 => n4640, IN3 => 
                           RAM_1_94_port, IN4 => n4629, IN5 => n4227, Q => 
                           n4230);
   U5538 : AO22X1 port map( IN1 => RAM_7_94_port, IN2 => n4662, IN3 => 
                           RAM_6_94_port, IN4 => n4651, Q => n4228);
   U5539 : AO221X1 port map( IN1 => RAM_4_94_port, IN2 => n4684, IN3 => 
                           RAM_5_94_port, IN4 => n4673, IN5 => n4228, Q => 
                           n4229);
   U5540 : OR4X1 port map( IN1 => n4232, IN2 => n4231, IN3 => n4230, IN4 => 
                           n4229, Q => RAMDOUT2(94));
   U5541 : AO22X1 port map( IN1 => RAM_11_95_port, IN2 => n4530, IN3 => 
                           RAM_10_95_port, IN4 => n4519, Q => n4233);
   U5542 : AO221X1 port map( IN1 => RAM_8_95_port, IN2 => n4552, IN3 => 
                           RAM_9_95_port, IN4 => n4541, IN5 => n4233, Q => 
                           n4240);
   U5543 : AO22X1 port map( IN1 => RAM_15_95_port, IN2 => n4574, IN3 => 
                           RAM_14_95_port, IN4 => n4563, Q => n4234);
   U5544 : AO221X1 port map( IN1 => RAM_12_95_port, IN2 => n4596, IN3 => 
                           RAM_13_95_port, IN4 => n4585, IN5 => n4234, Q => 
                           n4239);
   U5545 : AO22X1 port map( IN1 => RAM_3_95_port, IN2 => n4618, IN3 => 
                           RAM_2_95_port, IN4 => n4607, Q => n4235);
   U5546 : AO221X1 port map( IN1 => RAM_0_95_port, IN2 => n4640, IN3 => 
                           RAM_1_95_port, IN4 => n4629, IN5 => n4235, Q => 
                           n4238);
   U5547 : AO22X1 port map( IN1 => RAM_7_95_port, IN2 => n4662, IN3 => 
                           RAM_6_95_port, IN4 => n4651, Q => n4236);
   U5548 : AO221X1 port map( IN1 => RAM_4_95_port, IN2 => n4684, IN3 => 
                           RAM_5_95_port, IN4 => n4673, IN5 => n4236, Q => 
                           n4237);
   U5549 : AO22X1 port map( IN1 => RAM_11_96_port, IN2 => n4529, IN3 => 
                           RAM_10_96_port, IN4 => n4518, Q => n4241);
   U5550 : AO221X1 port map( IN1 => RAM_8_96_port, IN2 => n4551, IN3 => 
                           RAM_9_96_port, IN4 => n4540, IN5 => n4241, Q => 
                           n4248);
   U5551 : AO22X1 port map( IN1 => RAM_15_96_port, IN2 => n4573, IN3 => 
                           RAM_14_96_port, IN4 => n4562, Q => n4242);
   U5552 : AO221X1 port map( IN1 => RAM_12_96_port, IN2 => n4595, IN3 => 
                           RAM_13_96_port, IN4 => n4584, IN5 => n4242, Q => 
                           n4247);
   U5553 : AO22X1 port map( IN1 => RAM_3_96_port, IN2 => n4617, IN3 => 
                           RAM_2_96_port, IN4 => n4606, Q => n4243);
   U5554 : AO221X1 port map( IN1 => RAM_0_96_port, IN2 => n4639, IN3 => 
                           RAM_1_96_port, IN4 => n4628, IN5 => n4243, Q => 
                           n4246);
   U5555 : AO22X1 port map( IN1 => RAM_7_96_port, IN2 => n4661, IN3 => 
                           RAM_6_96_port, IN4 => n4650, Q => n4244);
   U5556 : AO221X1 port map( IN1 => RAM_4_96_port, IN2 => n4683, IN3 => 
                           RAM_5_96_port, IN4 => n4672, IN5 => n4244, Q => 
                           n4245);
   U5557 : OR4X1 port map( IN1 => n4248, IN2 => n4247, IN3 => n4246, IN4 => 
                           n4245, Q => RAMDOUT2(96));
   U5558 : AO22X1 port map( IN1 => RAM_11_97_port, IN2 => n4529, IN3 => 
                           RAM_10_97_port, IN4 => n4518, Q => n4249);
   U5559 : AO221X1 port map( IN1 => RAM_8_97_port, IN2 => n4551, IN3 => 
                           RAM_9_97_port, IN4 => n4540, IN5 => n4249, Q => 
                           n4256);
   U5560 : AO22X1 port map( IN1 => RAM_15_97_port, IN2 => n4573, IN3 => 
                           RAM_14_97_port, IN4 => n4562, Q => n4250);
   U5561 : AO221X1 port map( IN1 => RAM_12_97_port, IN2 => n4595, IN3 => 
                           RAM_13_97_port, IN4 => n4584, IN5 => n4250, Q => 
                           n4255);
   U5562 : AO22X1 port map( IN1 => RAM_3_97_port, IN2 => n4617, IN3 => 
                           RAM_2_97_port, IN4 => n4606, Q => n4251);
   U5563 : AO221X1 port map( IN1 => RAM_0_97_port, IN2 => n4639, IN3 => 
                           RAM_1_97_port, IN4 => n4628, IN5 => n4251, Q => 
                           n4254);
   U5564 : AO22X1 port map( IN1 => RAM_7_97_port, IN2 => n4661, IN3 => 
                           RAM_6_97_port, IN4 => n4650, Q => n4252);
   U5565 : AO221X1 port map( IN1 => RAM_4_97_port, IN2 => n4683, IN3 => 
                           RAM_5_97_port, IN4 => n4672, IN5 => n4252, Q => 
                           n4253);
   U5566 : OR4X1 port map( IN1 => n4256, IN2 => n4255, IN3 => n4254, IN4 => 
                           n4253, Q => RAMDOUT2(97));
   U5567 : AO22X1 port map( IN1 => RAM_11_98_port, IN2 => n4529, IN3 => 
                           RAM_10_98_port, IN4 => n4518, Q => n4257);
   U5568 : AO221X1 port map( IN1 => RAM_8_98_port, IN2 => n4551, IN3 => 
                           RAM_9_98_port, IN4 => n4540, IN5 => n4257, Q => 
                           n4264);
   U5569 : AO22X1 port map( IN1 => RAM_15_98_port, IN2 => n4573, IN3 => 
                           RAM_14_98_port, IN4 => n4562, Q => n4258);
   U5570 : AO221X1 port map( IN1 => RAM_12_98_port, IN2 => n4595, IN3 => 
                           RAM_13_98_port, IN4 => n4584, IN5 => n4258, Q => 
                           n4263);
   U5571 : AO22X1 port map( IN1 => RAM_3_98_port, IN2 => n4617, IN3 => 
                           RAM_2_98_port, IN4 => n4606, Q => n4259);
   U5572 : AO221X1 port map( IN1 => RAM_0_98_port, IN2 => n4639, IN3 => 
                           RAM_1_98_port, IN4 => n4628, IN5 => n4259, Q => 
                           n4262);
   U5573 : AO22X1 port map( IN1 => RAM_7_98_port, IN2 => n4661, IN3 => 
                           RAM_6_98_port, IN4 => n4650, Q => n4260);
   U5574 : AO221X1 port map( IN1 => RAM_4_98_port, IN2 => n4683, IN3 => 
                           RAM_5_98_port, IN4 => n4672, IN5 => n4260, Q => 
                           n4261);
   U5575 : OR4X1 port map( IN1 => n4264, IN2 => n4263, IN3 => n4262, IN4 => 
                           n4261, Q => RAMDOUT2(98));
   U5576 : AO22X1 port map( IN1 => RAM_11_99_port, IN2 => n4529, IN3 => 
                           RAM_10_99_port, IN4 => n4518, Q => n4265);
   U5577 : AO221X1 port map( IN1 => RAM_8_99_port, IN2 => n4551, IN3 => 
                           RAM_9_99_port, IN4 => n4540, IN5 => n4265, Q => 
                           n4272);
   U5578 : AO22X1 port map( IN1 => RAM_15_99_port, IN2 => n4573, IN3 => 
                           RAM_14_99_port, IN4 => n4562, Q => n4266);
   U5579 : AO221X1 port map( IN1 => RAM_12_99_port, IN2 => n4595, IN3 => 
                           RAM_13_99_port, IN4 => n4584, IN5 => n4266, Q => 
                           n4271);
   U5580 : AO22X1 port map( IN1 => RAM_3_99_port, IN2 => n4617, IN3 => 
                           RAM_2_99_port, IN4 => n4606, Q => n4267);
   U5581 : AO221X1 port map( IN1 => RAM_0_99_port, IN2 => n4639, IN3 => 
                           RAM_1_99_port, IN4 => n4628, IN5 => n4267, Q => 
                           n4270);
   U5582 : AO22X1 port map( IN1 => RAM_7_99_port, IN2 => n4661, IN3 => 
                           RAM_6_99_port, IN4 => n4650, Q => n4268);
   U5583 : AO221X1 port map( IN1 => RAM_4_99_port, IN2 => n4683, IN3 => 
                           RAM_5_99_port, IN4 => n4672, IN5 => n4268, Q => 
                           n4269);
   U5584 : OR4X1 port map( IN1 => n4272, IN2 => n4271, IN3 => n4270, IN4 => 
                           n4269, Q => RAMDOUT2(99));
   U5585 : AO22X1 port map( IN1 => RAM_11_100_port, IN2 => n4529, IN3 => 
                           RAM_10_100_port, IN4 => n4518, Q => n4273);
   U5586 : AO221X1 port map( IN1 => RAM_8_100_port, IN2 => n4551, IN3 => 
                           RAM_9_100_port, IN4 => n4540, IN5 => n4273, Q => 
                           n4280);
   U5587 : AO22X1 port map( IN1 => RAM_15_100_port, IN2 => n4573, IN3 => 
                           RAM_14_100_port, IN4 => n4562, Q => n4274);
   U5588 : AO221X1 port map( IN1 => RAM_12_100_port, IN2 => n4595, IN3 => 
                           RAM_13_100_port, IN4 => n4584, IN5 => n4274, Q => 
                           n4279);
   U5589 : AO22X1 port map( IN1 => RAM_3_100_port, IN2 => n4617, IN3 => 
                           RAM_2_100_port, IN4 => n4606, Q => n4275);
   U5590 : AO221X1 port map( IN1 => RAM_0_100_port, IN2 => n4639, IN3 => 
                           RAM_1_100_port, IN4 => n4628, IN5 => n4275, Q => 
                           n4278);
   U5591 : AO22X1 port map( IN1 => RAM_7_100_port, IN2 => n4661, IN3 => 
                           RAM_6_100_port, IN4 => n4650, Q => n4276);
   U5592 : AO221X1 port map( IN1 => RAM_4_100_port, IN2 => n4683, IN3 => 
                           RAM_5_100_port, IN4 => n4672, IN5 => n4276, Q => 
                           n4277);
   U5593 : OR4X1 port map( IN1 => n4280, IN2 => n4279, IN3 => n4278, IN4 => 
                           n4277, Q => RAMDOUT2(100));
   U5594 : AO22X1 port map( IN1 => RAM_11_101_port, IN2 => n4529, IN3 => 
                           RAM_10_101_port, IN4 => n4518, Q => n4281);
   U5595 : AO221X1 port map( IN1 => RAM_8_101_port, IN2 => n4551, IN3 => 
                           RAM_9_101_port, IN4 => n4540, IN5 => n4281, Q => 
                           n4288);
   U5596 : AO22X1 port map( IN1 => RAM_15_101_port, IN2 => n4573, IN3 => 
                           RAM_14_101_port, IN4 => n4562, Q => n4282);
   U5597 : AO221X1 port map( IN1 => RAM_12_101_port, IN2 => n4595, IN3 => 
                           RAM_13_101_port, IN4 => n4584, IN5 => n4282, Q => 
                           n4287);
   U5598 : AO22X1 port map( IN1 => RAM_3_101_port, IN2 => n4617, IN3 => 
                           RAM_2_101_port, IN4 => n4606, Q => n4283);
   U5599 : AO221X1 port map( IN1 => RAM_0_101_port, IN2 => n4639, IN3 => 
                           RAM_1_101_port, IN4 => n4628, IN5 => n4283, Q => 
                           n4286);
   U5600 : AO22X1 port map( IN1 => RAM_7_101_port, IN2 => n4661, IN3 => 
                           RAM_6_101_port, IN4 => n4650, Q => n4284);
   U5601 : AO221X1 port map( IN1 => RAM_4_101_port, IN2 => n4683, IN3 => 
                           RAM_5_101_port, IN4 => n4672, IN5 => n4284, Q => 
                           n4285);
   U5602 : OR4X1 port map( IN1 => n4288, IN2 => n4287, IN3 => n4286, IN4 => 
                           n4285, Q => RAMDOUT2(101));
   U5603 : AO22X1 port map( IN1 => RAM_11_102_port, IN2 => n4529, IN3 => 
                           RAM_10_102_port, IN4 => n4518, Q => n4289);
   U5604 : AO221X1 port map( IN1 => RAM_8_102_port, IN2 => n4551, IN3 => 
                           RAM_9_102_port, IN4 => n4540, IN5 => n4289, Q => 
                           n4296);
   U5605 : AO22X1 port map( IN1 => RAM_15_102_port, IN2 => n4573, IN3 => 
                           RAM_14_102_port, IN4 => n4562, Q => n4290);
   U5606 : AO221X1 port map( IN1 => RAM_12_102_port, IN2 => n4595, IN3 => 
                           RAM_13_102_port, IN4 => n4584, IN5 => n4290, Q => 
                           n4295);
   U5607 : AO22X1 port map( IN1 => RAM_3_102_port, IN2 => n4617, IN3 => 
                           RAM_2_102_port, IN4 => n4606, Q => n4291);
   U5608 : AO221X1 port map( IN1 => RAM_0_102_port, IN2 => n4639, IN3 => 
                           RAM_1_102_port, IN4 => n4628, IN5 => n4291, Q => 
                           n4294);
   U5609 : AO22X1 port map( IN1 => RAM_7_102_port, IN2 => n4661, IN3 => 
                           RAM_6_102_port, IN4 => n4650, Q => n4292);
   U5610 : AO221X1 port map( IN1 => RAM_4_102_port, IN2 => n4683, IN3 => 
                           RAM_5_102_port, IN4 => n4672, IN5 => n4292, Q => 
                           n4293);
   U5611 : OR4X1 port map( IN1 => n4296, IN2 => n4295, IN3 => n4294, IN4 => 
                           n4293, Q => RAMDOUT2(102));
   U5612 : AO22X1 port map( IN1 => RAM_11_103_port, IN2 => n4529, IN3 => 
                           RAM_10_103_port, IN4 => n4518, Q => n4297);
   U5613 : AO221X1 port map( IN1 => RAM_8_103_port, IN2 => n4551, IN3 => 
                           RAM_9_103_port, IN4 => n4540, IN5 => n4297, Q => 
                           n4304);
   U5614 : AO22X1 port map( IN1 => RAM_15_103_port, IN2 => n4573, IN3 => 
                           RAM_14_103_port, IN4 => n4562, Q => n4298);
   U5615 : AO221X1 port map( IN1 => RAM_12_103_port, IN2 => n4595, IN3 => 
                           RAM_13_103_port, IN4 => n4584, IN5 => n4298, Q => 
                           n4303);
   U5616 : AO22X1 port map( IN1 => RAM_3_103_port, IN2 => n4617, IN3 => 
                           RAM_2_103_port, IN4 => n4606, Q => n4299);
   U5617 : AO221X1 port map( IN1 => RAM_0_103_port, IN2 => n4639, IN3 => 
                           RAM_1_103_port, IN4 => n4628, IN5 => n4299, Q => 
                           n4302);
   U5618 : AO22X1 port map( IN1 => RAM_7_103_port, IN2 => n4661, IN3 => 
                           RAM_6_103_port, IN4 => n4650, Q => n4300);
   U5619 : AO221X1 port map( IN1 => RAM_4_103_port, IN2 => n4683, IN3 => 
                           RAM_5_103_port, IN4 => n4672, IN5 => n4300, Q => 
                           n4301);
   U5620 : OR4X1 port map( IN1 => n4304, IN2 => n4303, IN3 => n4302, IN4 => 
                           n4301, Q => RAMDOUT2(103));
   U5621 : AO22X1 port map( IN1 => RAM_11_104_port, IN2 => n4529, IN3 => 
                           RAM_10_104_port, IN4 => n4518, Q => n4305);
   U5622 : AO221X1 port map( IN1 => RAM_8_104_port, IN2 => n4551, IN3 => 
                           RAM_9_104_port, IN4 => n4540, IN5 => n4305, Q => 
                           n4312);
   U5623 : AO22X1 port map( IN1 => RAM_15_104_port, IN2 => n4573, IN3 => 
                           RAM_14_104_port, IN4 => n4562, Q => n4306);
   U5624 : AO221X1 port map( IN1 => RAM_12_104_port, IN2 => n4595, IN3 => 
                           RAM_13_104_port, IN4 => n4584, IN5 => n4306, Q => 
                           n4311);
   U5625 : AO22X1 port map( IN1 => RAM_3_104_port, IN2 => n4617, IN3 => 
                           RAM_2_104_port, IN4 => n4606, Q => n4307);
   U5626 : AO221X1 port map( IN1 => RAM_0_104_port, IN2 => n4639, IN3 => 
                           RAM_1_104_port, IN4 => n4628, IN5 => n4307, Q => 
                           n4310);
   U5627 : AO22X1 port map( IN1 => RAM_7_104_port, IN2 => n4661, IN3 => 
                           RAM_6_104_port, IN4 => n4650, Q => n4308);
   U5628 : AO221X1 port map( IN1 => RAM_4_104_port, IN2 => n4683, IN3 => 
                           RAM_5_104_port, IN4 => n4672, IN5 => n4308, Q => 
                           n4309);
   U5629 : OR4X1 port map( IN1 => n4312, IN2 => n4311, IN3 => n4310, IN4 => 
                           n4309, Q => RAMDOUT2(104));
   U5630 : AO22X1 port map( IN1 => RAM_11_105_port, IN2 => n4529, IN3 => 
                           RAM_10_105_port, IN4 => n4518, Q => n4313);
   U5631 : AO221X1 port map( IN1 => RAM_8_105_port, IN2 => n4551, IN3 => 
                           RAM_9_105_port, IN4 => n4540, IN5 => n4313, Q => 
                           n4320);
   U5632 : AO22X1 port map( IN1 => RAM_15_105_port, IN2 => n4573, IN3 => 
                           RAM_14_105_port, IN4 => n4562, Q => n4314);
   U5633 : AO221X1 port map( IN1 => RAM_12_105_port, IN2 => n4595, IN3 => 
                           RAM_13_105_port, IN4 => n4584, IN5 => n4314, Q => 
                           n4319);
   U5634 : AO22X1 port map( IN1 => RAM_3_105_port, IN2 => n4617, IN3 => 
                           RAM_2_105_port, IN4 => n4606, Q => n4315);
   U5635 : AO221X1 port map( IN1 => RAM_0_105_port, IN2 => n4639, IN3 => 
                           RAM_1_105_port, IN4 => n4628, IN5 => n4315, Q => 
                           n4318);
   U5636 : AO22X1 port map( IN1 => RAM_7_105_port, IN2 => n4661, IN3 => 
                           RAM_6_105_port, IN4 => n4650, Q => n4316);
   U5637 : AO221X1 port map( IN1 => RAM_4_105_port, IN2 => n4683, IN3 => 
                           RAM_5_105_port, IN4 => n4672, IN5 => n4316, Q => 
                           n4317);
   U5638 : OR4X1 port map( IN1 => n4320, IN2 => n4319, IN3 => n4318, IN4 => 
                           n4317, Q => RAMDOUT2(105));
   U5639 : AO22X1 port map( IN1 => RAM_11_106_port, IN2 => n4529, IN3 => 
                           RAM_10_106_port, IN4 => n4518, Q => n4321);
   U5640 : AO221X1 port map( IN1 => RAM_8_106_port, IN2 => n4551, IN3 => 
                           RAM_9_106_port, IN4 => n4540, IN5 => n4321, Q => 
                           n4328);
   U5641 : AO22X1 port map( IN1 => RAM_15_106_port, IN2 => n4573, IN3 => 
                           RAM_14_106_port, IN4 => n4562, Q => n4322);
   U5642 : AO221X1 port map( IN1 => RAM_12_106_port, IN2 => n4595, IN3 => 
                           RAM_13_106_port, IN4 => n4584, IN5 => n4322, Q => 
                           n4327);
   U5643 : AO22X1 port map( IN1 => RAM_3_106_port, IN2 => n4617, IN3 => 
                           RAM_2_106_port, IN4 => n4606, Q => n4323);
   U5644 : AO221X1 port map( IN1 => RAM_0_106_port, IN2 => n4639, IN3 => 
                           RAM_1_106_port, IN4 => n4628, IN5 => n4323, Q => 
                           n4326);
   U5645 : AO22X1 port map( IN1 => RAM_7_106_port, IN2 => n4661, IN3 => 
                           RAM_6_106_port, IN4 => n4650, Q => n4324);
   U5646 : AO221X1 port map( IN1 => RAM_4_106_port, IN2 => n4683, IN3 => 
                           RAM_5_106_port, IN4 => n4672, IN5 => n4324, Q => 
                           n4325);
   U5647 : OR4X1 port map( IN1 => n4328, IN2 => n4327, IN3 => n4326, IN4 => 
                           n4325, Q => RAMDOUT2(106));
   U5648 : AO22X1 port map( IN1 => RAM_11_107_port, IN2 => n4529, IN3 => 
                           RAM_10_107_port, IN4 => n4518, Q => n4329);
   U5649 : AO221X1 port map( IN1 => RAM_8_107_port, IN2 => n4551, IN3 => 
                           RAM_9_107_port, IN4 => n4540, IN5 => n4329, Q => 
                           n4336);
   U5650 : AO22X1 port map( IN1 => RAM_15_107_port, IN2 => n4573, IN3 => 
                           RAM_14_107_port, IN4 => n4562, Q => n4330);
   U5651 : AO221X1 port map( IN1 => RAM_12_107_port, IN2 => n4595, IN3 => 
                           RAM_13_107_port, IN4 => n4584, IN5 => n4330, Q => 
                           n4335);
   U5652 : AO22X1 port map( IN1 => RAM_3_107_port, IN2 => n4617, IN3 => 
                           RAM_2_107_port, IN4 => n4606, Q => n4331);
   U5653 : AO221X1 port map( IN1 => RAM_0_107_port, IN2 => n4639, IN3 => 
                           RAM_1_107_port, IN4 => n4628, IN5 => n4331, Q => 
                           n4334);
   U5654 : AO22X1 port map( IN1 => RAM_7_107_port, IN2 => n4661, IN3 => 
                           RAM_6_107_port, IN4 => n4650, Q => n4332);
   U5655 : AO221X1 port map( IN1 => RAM_4_107_port, IN2 => n4683, IN3 => 
                           RAM_5_107_port, IN4 => n4672, IN5 => n4332, Q => 
                           n4333);
   U5656 : OR4X1 port map( IN1 => n4336, IN2 => n4335, IN3 => n4334, IN4 => 
                           n4333, Q => RAMDOUT2(107));
   U5657 : AO22X1 port map( IN1 => RAM_11_108_port, IN2 => n4528, IN3 => 
                           RAM_10_108_port, IN4 => n4517, Q => n4337);
   U5658 : AO221X1 port map( IN1 => RAM_8_108_port, IN2 => n4550, IN3 => 
                           RAM_9_108_port, IN4 => n4539, IN5 => n4337, Q => 
                           n4344);
   U5659 : AO22X1 port map( IN1 => RAM_15_108_port, IN2 => n4572, IN3 => 
                           RAM_14_108_port, IN4 => n4561, Q => n4338);
   U5660 : AO221X1 port map( IN1 => RAM_12_108_port, IN2 => n4594, IN3 => 
                           RAM_13_108_port, IN4 => n4583, IN5 => n4338, Q => 
                           n4343);
   U5661 : AO22X1 port map( IN1 => RAM_3_108_port, IN2 => n4616, IN3 => 
                           RAM_2_108_port, IN4 => n4605, Q => n4339);
   U5662 : AO221X1 port map( IN1 => RAM_0_108_port, IN2 => n4638, IN3 => 
                           RAM_1_108_port, IN4 => n4627, IN5 => n4339, Q => 
                           n4342);
   U5663 : AO22X1 port map( IN1 => RAM_7_108_port, IN2 => n4660, IN3 => 
                           RAM_6_108_port, IN4 => n4649, Q => n4340);
   U5664 : AO221X1 port map( IN1 => RAM_4_108_port, IN2 => n4682, IN3 => 
                           RAM_5_108_port, IN4 => n4671, IN5 => n4340, Q => 
                           n4341);
   U5665 : OR4X1 port map( IN1 => n4344, IN2 => n4343, IN3 => n4342, IN4 => 
                           n4341, Q => RAMDOUT2(108));
   U5666 : AO22X1 port map( IN1 => RAM_11_109_port, IN2 => n4528, IN3 => 
                           RAM_10_109_port, IN4 => n4517, Q => n4345);
   U5667 : AO221X1 port map( IN1 => RAM_8_109_port, IN2 => n4550, IN3 => 
                           RAM_9_109_port, IN4 => n4539, IN5 => n4345, Q => 
                           n4352);
   U5668 : AO22X1 port map( IN1 => RAM_15_109_port, IN2 => n4572, IN3 => 
                           RAM_14_109_port, IN4 => n4561, Q => n4346);
   U5669 : AO221X1 port map( IN1 => RAM_12_109_port, IN2 => n4594, IN3 => 
                           RAM_13_109_port, IN4 => n4583, IN5 => n4346, Q => 
                           n4351);
   U5670 : AO22X1 port map( IN1 => RAM_3_109_port, IN2 => n4616, IN3 => 
                           RAM_2_109_port, IN4 => n4605, Q => n4347);
   U5671 : AO221X1 port map( IN1 => RAM_0_109_port, IN2 => n4638, IN3 => 
                           RAM_1_109_port, IN4 => n4627, IN5 => n4347, Q => 
                           n4350);
   U5672 : AO22X1 port map( IN1 => RAM_7_109_port, IN2 => n4660, IN3 => 
                           RAM_6_109_port, IN4 => n4649, Q => n4348);
   U5673 : AO221X1 port map( IN1 => RAM_4_109_port, IN2 => n4682, IN3 => 
                           RAM_5_109_port, IN4 => n4671, IN5 => n4348, Q => 
                           n4349);
   U5674 : OR4X1 port map( IN1 => n4352, IN2 => n4351, IN3 => n4350, IN4 => 
                           n4349, Q => RAMDOUT2(109));
   U5675 : AO22X1 port map( IN1 => RAM_11_110_port, IN2 => n4528, IN3 => 
                           RAM_10_110_port, IN4 => n4517, Q => n4353);
   U5676 : AO221X1 port map( IN1 => RAM_8_110_port, IN2 => n4550, IN3 => 
                           RAM_9_110_port, IN4 => n4539, IN5 => n4353, Q => 
                           n4360);
   U5677 : AO22X1 port map( IN1 => RAM_15_110_port, IN2 => n4572, IN3 => 
                           RAM_14_110_port, IN4 => n4561, Q => n4354);
   U5678 : AO221X1 port map( IN1 => RAM_12_110_port, IN2 => n4594, IN3 => 
                           RAM_13_110_port, IN4 => n4583, IN5 => n4354, Q => 
                           n4359);
   U5679 : AO22X1 port map( IN1 => RAM_3_110_port, IN2 => n4616, IN3 => 
                           RAM_2_110_port, IN4 => n4605, Q => n4355);
   U5680 : AO221X1 port map( IN1 => RAM_0_110_port, IN2 => n4638, IN3 => 
                           RAM_1_110_port, IN4 => n4627, IN5 => n4355, Q => 
                           n4358);
   U5681 : AO22X1 port map( IN1 => RAM_7_110_port, IN2 => n4660, IN3 => 
                           RAM_6_110_port, IN4 => n4649, Q => n4356);
   U5682 : AO221X1 port map( IN1 => RAM_4_110_port, IN2 => n4682, IN3 => 
                           RAM_5_110_port, IN4 => n4671, IN5 => n4356, Q => 
                           n4357);
   U5683 : OR4X1 port map( IN1 => n4360, IN2 => n4359, IN3 => n4358, IN4 => 
                           n4357, Q => RAMDOUT2(110));
   U5684 : AO22X1 port map( IN1 => RAM_11_111_port, IN2 => n4528, IN3 => 
                           RAM_10_111_port, IN4 => n4517, Q => n4361);
   U5685 : AO221X1 port map( IN1 => RAM_8_111_port, IN2 => n4550, IN3 => 
                           RAM_9_111_port, IN4 => n4539, IN5 => n4361, Q => 
                           n4368);
   U5686 : AO22X1 port map( IN1 => RAM_15_111_port, IN2 => n4572, IN3 => 
                           RAM_14_111_port, IN4 => n4561, Q => n4362);
   U5687 : AO221X1 port map( IN1 => RAM_12_111_port, IN2 => n4594, IN3 => 
                           RAM_13_111_port, IN4 => n4583, IN5 => n4362, Q => 
                           n4367);
   U5688 : AO22X1 port map( IN1 => RAM_3_111_port, IN2 => n4616, IN3 => 
                           RAM_2_111_port, IN4 => n4605, Q => n4363);
   U5689 : AO221X1 port map( IN1 => RAM_0_111_port, IN2 => n4638, IN3 => 
                           RAM_1_111_port, IN4 => n4627, IN5 => n4363, Q => 
                           n4366);
   U5690 : AO22X1 port map( IN1 => RAM_7_111_port, IN2 => n4660, IN3 => 
                           RAM_6_111_port, IN4 => n4649, Q => n4364);
   U5691 : AO221X1 port map( IN1 => RAM_4_111_port, IN2 => n4682, IN3 => 
                           RAM_5_111_port, IN4 => n4671, IN5 => n4364, Q => 
                           n4365);
   U5692 : OR4X1 port map( IN1 => n4368, IN2 => n4367, IN3 => n4366, IN4 => 
                           n4365, Q => RAMDOUT2(111));
   U5693 : AO22X1 port map( IN1 => RAM_11_112_port, IN2 => n4528, IN3 => 
                           RAM_10_112_port, IN4 => n4517, Q => n4369);
   U5694 : AO221X1 port map( IN1 => RAM_8_112_port, IN2 => n4550, IN3 => 
                           RAM_9_112_port, IN4 => n4539, IN5 => n4369, Q => 
                           n4376);
   U5695 : AO22X1 port map( IN1 => RAM_15_112_port, IN2 => n4572, IN3 => 
                           RAM_14_112_port, IN4 => n4561, Q => n4370);
   U5696 : AO221X1 port map( IN1 => RAM_12_112_port, IN2 => n4594, IN3 => 
                           RAM_13_112_port, IN4 => n4583, IN5 => n4370, Q => 
                           n4375);
   U5697 : AO22X1 port map( IN1 => RAM_3_112_port, IN2 => n4616, IN3 => 
                           RAM_2_112_port, IN4 => n4605, Q => n4371);
   U5698 : AO221X1 port map( IN1 => RAM_0_112_port, IN2 => n4638, IN3 => 
                           RAM_1_112_port, IN4 => n4627, IN5 => n4371, Q => 
                           n4374);
   U5699 : AO22X1 port map( IN1 => RAM_7_112_port, IN2 => n4660, IN3 => 
                           RAM_6_112_port, IN4 => n4649, Q => n4372);
   U5700 : AO221X1 port map( IN1 => RAM_4_112_port, IN2 => n4682, IN3 => 
                           RAM_5_112_port, IN4 => n4671, IN5 => n4372, Q => 
                           n4373);
   U5701 : OR4X1 port map( IN1 => n4376, IN2 => n4375, IN3 => n4374, IN4 => 
                           n4373, Q => RAMDOUT2(112));
   U5702 : AO22X1 port map( IN1 => RAM_11_113_port, IN2 => n4528, IN3 => 
                           RAM_10_113_port, IN4 => n4517, Q => n4377);
   U5703 : AO221X1 port map( IN1 => RAM_8_113_port, IN2 => n4550, IN3 => 
                           RAM_9_113_port, IN4 => n4539, IN5 => n4377, Q => 
                           n4384);
   U5704 : AO22X1 port map( IN1 => RAM_15_113_port, IN2 => n4572, IN3 => 
                           RAM_14_113_port, IN4 => n4561, Q => n4378);
   U5705 : AO221X1 port map( IN1 => RAM_12_113_port, IN2 => n4594, IN3 => 
                           RAM_13_113_port, IN4 => n4583, IN5 => n4378, Q => 
                           n4383);
   U5706 : AO22X1 port map( IN1 => RAM_3_113_port, IN2 => n4616, IN3 => 
                           RAM_2_113_port, IN4 => n4605, Q => n4379);
   U5707 : AO221X1 port map( IN1 => RAM_0_113_port, IN2 => n4638, IN3 => 
                           RAM_1_113_port, IN4 => n4627, IN5 => n4379, Q => 
                           n4382);
   U5708 : AO22X1 port map( IN1 => RAM_7_113_port, IN2 => n4660, IN3 => 
                           RAM_6_113_port, IN4 => n4649, Q => n4380);
   U5709 : AO221X1 port map( IN1 => RAM_4_113_port, IN2 => n4682, IN3 => 
                           RAM_5_113_port, IN4 => n4671, IN5 => n4380, Q => 
                           n4381);
   U5710 : OR4X1 port map( IN1 => n4384, IN2 => n4383, IN3 => n4382, IN4 => 
                           n4381, Q => RAMDOUT2(113));
   U5711 : AO22X1 port map( IN1 => RAM_11_114_port, IN2 => n4528, IN3 => 
                           RAM_10_114_port, IN4 => n4517, Q => n4385);
   U5712 : AO221X1 port map( IN1 => RAM_8_114_port, IN2 => n4550, IN3 => 
                           RAM_9_114_port, IN4 => n4539, IN5 => n4385, Q => 
                           n4392);
   U5713 : AO22X1 port map( IN1 => RAM_15_114_port, IN2 => n4572, IN3 => 
                           RAM_14_114_port, IN4 => n4561, Q => n4386);
   U5714 : AO221X1 port map( IN1 => RAM_12_114_port, IN2 => n4594, IN3 => 
                           RAM_13_114_port, IN4 => n4583, IN5 => n4386, Q => 
                           n4391);
   U5715 : AO22X1 port map( IN1 => RAM_3_114_port, IN2 => n4616, IN3 => 
                           RAM_2_114_port, IN4 => n4605, Q => n4387);
   U5716 : AO221X1 port map( IN1 => RAM_0_114_port, IN2 => n4638, IN3 => 
                           RAM_1_114_port, IN4 => n4627, IN5 => n4387, Q => 
                           n4390);
   U5717 : AO22X1 port map( IN1 => RAM_7_114_port, IN2 => n4660, IN3 => 
                           RAM_6_114_port, IN4 => n4649, Q => n4388);
   U5718 : AO221X1 port map( IN1 => RAM_4_114_port, IN2 => n4682, IN3 => 
                           RAM_5_114_port, IN4 => n4671, IN5 => n4388, Q => 
                           n4389);
   U5719 : OR4X1 port map( IN1 => n4392, IN2 => n4391, IN3 => n4390, IN4 => 
                           n4389, Q => RAMDOUT2(114));
   U5720 : AO22X1 port map( IN1 => RAM_11_115_port, IN2 => n4528, IN3 => 
                           RAM_10_115_port, IN4 => n4517, Q => n4393);
   U5721 : AO221X1 port map( IN1 => RAM_8_115_port, IN2 => n4550, IN3 => 
                           RAM_9_115_port, IN4 => n4539, IN5 => n4393, Q => 
                           n4400);
   U5722 : AO22X1 port map( IN1 => RAM_15_115_port, IN2 => n4572, IN3 => 
                           RAM_14_115_port, IN4 => n4561, Q => n4394);
   U5723 : AO221X1 port map( IN1 => RAM_12_115_port, IN2 => n4594, IN3 => 
                           RAM_13_115_port, IN4 => n4583, IN5 => n4394, Q => 
                           n4399);
   U5724 : AO22X1 port map( IN1 => RAM_3_115_port, IN2 => n4616, IN3 => 
                           RAM_2_115_port, IN4 => n4605, Q => n4395);
   U5725 : AO221X1 port map( IN1 => RAM_0_115_port, IN2 => n4638, IN3 => 
                           RAM_1_115_port, IN4 => n4627, IN5 => n4395, Q => 
                           n4398);
   U5726 : AO22X1 port map( IN1 => RAM_7_115_port, IN2 => n4660, IN3 => 
                           RAM_6_115_port, IN4 => n4649, Q => n4396);
   U5727 : AO221X1 port map( IN1 => RAM_4_115_port, IN2 => n4682, IN3 => 
                           RAM_5_115_port, IN4 => n4671, IN5 => n4396, Q => 
                           n4397);
   U5728 : OR4X1 port map( IN1 => n4400, IN2 => n4399, IN3 => n4398, IN4 => 
                           n4397, Q => RAMDOUT2(115));
   U5729 : AO22X1 port map( IN1 => RAM_11_116_port, IN2 => n4528, IN3 => 
                           RAM_10_116_port, IN4 => n4517, Q => n4401);
   U5730 : AO221X1 port map( IN1 => RAM_8_116_port, IN2 => n4550, IN3 => 
                           RAM_9_116_port, IN4 => n4539, IN5 => n4401, Q => 
                           n4408);
   U5731 : AO22X1 port map( IN1 => RAM_15_116_port, IN2 => n4572, IN3 => 
                           RAM_14_116_port, IN4 => n4561, Q => n4402);
   U5732 : AO221X1 port map( IN1 => RAM_12_116_port, IN2 => n4594, IN3 => 
                           RAM_13_116_port, IN4 => n4583, IN5 => n4402, Q => 
                           n4407);
   U5733 : AO22X1 port map( IN1 => RAM_3_116_port, IN2 => n4616, IN3 => 
                           RAM_2_116_port, IN4 => n4605, Q => n4403);
   U5734 : AO221X1 port map( IN1 => RAM_0_116_port, IN2 => n4638, IN3 => 
                           RAM_1_116_port, IN4 => n4627, IN5 => n4403, Q => 
                           n4406);
   U5735 : AO22X1 port map( IN1 => RAM_7_116_port, IN2 => n4660, IN3 => 
                           RAM_6_116_port, IN4 => n4649, Q => n4404);
   U5736 : AO221X1 port map( IN1 => RAM_4_116_port, IN2 => n4682, IN3 => 
                           RAM_5_116_port, IN4 => n4671, IN5 => n4404, Q => 
                           n4405);
   U5737 : OR4X1 port map( IN1 => n4408, IN2 => n4407, IN3 => n4406, IN4 => 
                           n4405, Q => RAMDOUT2(116));
   U5738 : AO22X1 port map( IN1 => RAM_11_117_port, IN2 => n4528, IN3 => 
                           RAM_10_117_port, IN4 => n4517, Q => n4409);
   U5739 : AO221X1 port map( IN1 => RAM_8_117_port, IN2 => n4550, IN3 => 
                           RAM_9_117_port, IN4 => n4539, IN5 => n4409, Q => 
                           n4416);
   U5740 : AO22X1 port map( IN1 => RAM_15_117_port, IN2 => n4572, IN3 => 
                           RAM_14_117_port, IN4 => n4561, Q => n4410);
   U5741 : AO221X1 port map( IN1 => RAM_12_117_port, IN2 => n4594, IN3 => 
                           RAM_13_117_port, IN4 => n4583, IN5 => n4410, Q => 
                           n4415);
   U5742 : AO22X1 port map( IN1 => RAM_3_117_port, IN2 => n4616, IN3 => 
                           RAM_2_117_port, IN4 => n4605, Q => n4411);
   U5743 : AO221X1 port map( IN1 => RAM_0_117_port, IN2 => n4638, IN3 => 
                           RAM_1_117_port, IN4 => n4627, IN5 => n4411, Q => 
                           n4414);
   U5744 : AO22X1 port map( IN1 => RAM_7_117_port, IN2 => n4660, IN3 => 
                           RAM_6_117_port, IN4 => n4649, Q => n4412);
   U5745 : AO221X1 port map( IN1 => RAM_4_117_port, IN2 => n4682, IN3 => 
                           RAM_5_117_port, IN4 => n4671, IN5 => n4412, Q => 
                           n4413);
   U5746 : OR4X1 port map( IN1 => n4416, IN2 => n4415, IN3 => n4414, IN4 => 
                           n4413, Q => RAMDOUT2(117));
   U5747 : AO22X1 port map( IN1 => RAM_11_118_port, IN2 => n4528, IN3 => 
                           RAM_10_118_port, IN4 => n4517, Q => n4417);
   U5748 : AO221X1 port map( IN1 => RAM_8_118_port, IN2 => n4550, IN3 => 
                           RAM_9_118_port, IN4 => n4539, IN5 => n4417, Q => 
                           n4424);
   U5749 : AO22X1 port map( IN1 => RAM_15_118_port, IN2 => n4572, IN3 => 
                           RAM_14_118_port, IN4 => n4561, Q => n4418);
   U5750 : AO221X1 port map( IN1 => RAM_12_118_port, IN2 => n4594, IN3 => 
                           RAM_13_118_port, IN4 => n4583, IN5 => n4418, Q => 
                           n4423);
   U5751 : AO22X1 port map( IN1 => RAM_3_118_port, IN2 => n4616, IN3 => 
                           RAM_2_118_port, IN4 => n4605, Q => n4419);
   U5752 : AO221X1 port map( IN1 => RAM_0_118_port, IN2 => n4638, IN3 => 
                           RAM_1_118_port, IN4 => n4627, IN5 => n4419, Q => 
                           n4422);
   U5753 : AO22X1 port map( IN1 => RAM_7_118_port, IN2 => n4660, IN3 => 
                           RAM_6_118_port, IN4 => n4649, Q => n4420);
   U5754 : AO221X1 port map( IN1 => RAM_4_118_port, IN2 => n4682, IN3 => 
                           RAM_5_118_port, IN4 => n4671, IN5 => n4420, Q => 
                           n4421);
   U5755 : OR4X1 port map( IN1 => n4424, IN2 => n4423, IN3 => n4422, IN4 => 
                           n4421, Q => RAMDOUT2(118));
   U5756 : AO22X1 port map( IN1 => RAM_11_119_port, IN2 => n4528, IN3 => 
                           RAM_10_119_port, IN4 => n4517, Q => n4425);
   U5757 : AO221X1 port map( IN1 => RAM_8_119_port, IN2 => n4550, IN3 => 
                           RAM_9_119_port, IN4 => n4539, IN5 => n4425, Q => 
                           n4432);
   U5758 : AO22X1 port map( IN1 => RAM_15_119_port, IN2 => n4572, IN3 => 
                           RAM_14_119_port, IN4 => n4561, Q => n4426);
   U5759 : AO221X1 port map( IN1 => RAM_12_119_port, IN2 => n4594, IN3 => 
                           RAM_13_119_port, IN4 => n4583, IN5 => n4426, Q => 
                           n4431);
   U5760 : AO22X1 port map( IN1 => RAM_3_119_port, IN2 => n4616, IN3 => 
                           RAM_2_119_port, IN4 => n4605, Q => n4427);
   U5761 : AO221X1 port map( IN1 => RAM_0_119_port, IN2 => n4638, IN3 => 
                           RAM_1_119_port, IN4 => n4627, IN5 => n4427, Q => 
                           n4430);
   U5762 : AO22X1 port map( IN1 => RAM_7_119_port, IN2 => n4660, IN3 => 
                           RAM_6_119_port, IN4 => n4649, Q => n4428);
   U5763 : AO221X1 port map( IN1 => RAM_4_119_port, IN2 => n4682, IN3 => 
                           RAM_5_119_port, IN4 => n4671, IN5 => n4428, Q => 
                           n4429);
   U5764 : OR4X1 port map( IN1 => n4432, IN2 => n4431, IN3 => n4430, IN4 => 
                           n4429, Q => RAMDOUT2(119));
   U5765 : AO22X1 port map( IN1 => RAM_11_120_port, IN2 => n4527, IN3 => 
                           RAM_10_120_port, IN4 => n4516, Q => n4433);
   U5766 : AO221X1 port map( IN1 => RAM_8_120_port, IN2 => n4549, IN3 => 
                           RAM_9_120_port, IN4 => n4538, IN5 => n4433, Q => 
                           n4440);
   U5767 : AO22X1 port map( IN1 => RAM_15_120_port, IN2 => n4571, IN3 => 
                           RAM_14_120_port, IN4 => n4560, Q => n4434);
   U5768 : AO221X1 port map( IN1 => RAM_12_120_port, IN2 => n4593, IN3 => 
                           RAM_13_120_port, IN4 => n4582, IN5 => n4434, Q => 
                           n4439);
   U5769 : AO22X1 port map( IN1 => RAM_3_120_port, IN2 => n4615, IN3 => 
                           RAM_2_120_port, IN4 => n4604, Q => n4435);
   U5770 : AO221X1 port map( IN1 => RAM_0_120_port, IN2 => n4637, IN3 => 
                           RAM_1_120_port, IN4 => n4626, IN5 => n4435, Q => 
                           n4438);
   U5771 : AO22X1 port map( IN1 => RAM_7_120_port, IN2 => n4659, IN3 => 
                           RAM_6_120_port, IN4 => n4648, Q => n4436);
   U5772 : AO221X1 port map( IN1 => RAM_4_120_port, IN2 => n4681, IN3 => 
                           RAM_5_120_port, IN4 => n4670, IN5 => n4436, Q => 
                           n4437);
   U5773 : OR4X1 port map( IN1 => n4440, IN2 => n4439, IN3 => n4438, IN4 => 
                           n4437, Q => RAMDOUT2(120));
   U5774 : AO22X1 port map( IN1 => RAM_11_121_port, IN2 => n4527, IN3 => 
                           RAM_10_121_port, IN4 => n4516, Q => n4441);
   U5775 : AO221X1 port map( IN1 => RAM_8_121_port, IN2 => n4549, IN3 => 
                           RAM_9_121_port, IN4 => n4538, IN5 => n4441, Q => 
                           n4448);
   U5776 : AO22X1 port map( IN1 => RAM_15_121_port, IN2 => n4571, IN3 => 
                           RAM_14_121_port, IN4 => n4560, Q => n4442);
   U5777 : AO221X1 port map( IN1 => RAM_12_121_port, IN2 => n4593, IN3 => 
                           RAM_13_121_port, IN4 => n4582, IN5 => n4442, Q => 
                           n4447);
   U5778 : AO22X1 port map( IN1 => RAM_3_121_port, IN2 => n4615, IN3 => 
                           RAM_2_121_port, IN4 => n4604, Q => n4443);
   U5779 : AO221X1 port map( IN1 => RAM_0_121_port, IN2 => n4637, IN3 => 
                           RAM_1_121_port, IN4 => n4626, IN5 => n4443, Q => 
                           n4446);
   U5780 : AO22X1 port map( IN1 => RAM_7_121_port, IN2 => n4659, IN3 => 
                           RAM_6_121_port, IN4 => n4648, Q => n4444);
   U5781 : AO221X1 port map( IN1 => RAM_4_121_port, IN2 => n4681, IN3 => 
                           RAM_5_121_port, IN4 => n4670, IN5 => n4444, Q => 
                           n4445);
   U5782 : OR4X1 port map( IN1 => n4448, IN2 => n4447, IN3 => n4446, IN4 => 
                           n4445, Q => RAMDOUT2(121));
   U5783 : AO22X1 port map( IN1 => RAM_11_122_port, IN2 => n4527, IN3 => 
                           RAM_10_122_port, IN4 => n4516, Q => n4449);
   U5784 : AO221X1 port map( IN1 => RAM_8_122_port, IN2 => n4549, IN3 => 
                           RAM_9_122_port, IN4 => n4538, IN5 => n4449, Q => 
                           n4456);
   U5785 : AO22X1 port map( IN1 => RAM_15_122_port, IN2 => n4571, IN3 => 
                           RAM_14_122_port, IN4 => n4560, Q => n4450);
   U5786 : AO221X1 port map( IN1 => RAM_12_122_port, IN2 => n4593, IN3 => 
                           RAM_13_122_port, IN4 => n4582, IN5 => n4450, Q => 
                           n4455);
   U5787 : AO22X1 port map( IN1 => RAM_3_122_port, IN2 => n4615, IN3 => 
                           RAM_2_122_port, IN4 => n4604, Q => n4451);
   U5788 : AO221X1 port map( IN1 => RAM_0_122_port, IN2 => n4637, IN3 => 
                           RAM_1_122_port, IN4 => n4626, IN5 => n4451, Q => 
                           n4454);
   U5789 : AO22X1 port map( IN1 => RAM_7_122_port, IN2 => n4659, IN3 => 
                           RAM_6_122_port, IN4 => n4648, Q => n4452);
   U5790 : AO221X1 port map( IN1 => RAM_4_122_port, IN2 => n4681, IN3 => 
                           RAM_5_122_port, IN4 => n4670, IN5 => n4452, Q => 
                           n4453);
   U5791 : OR4X1 port map( IN1 => n4456, IN2 => n4455, IN3 => n4454, IN4 => 
                           n4453, Q => RAMDOUT2(122));
   U5792 : AO22X1 port map( IN1 => RAM_11_123_port, IN2 => n4527, IN3 => 
                           RAM_10_123_port, IN4 => n4516, Q => n4457);
   U5793 : AO221X1 port map( IN1 => RAM_8_123_port, IN2 => n4549, IN3 => 
                           RAM_9_123_port, IN4 => n4538, IN5 => n4457, Q => 
                           n4464);
   U5794 : AO22X1 port map( IN1 => RAM_15_123_port, IN2 => n4571, IN3 => 
                           RAM_14_123_port, IN4 => n4560, Q => n4458);
   U5795 : AO221X1 port map( IN1 => RAM_12_123_port, IN2 => n4593, IN3 => 
                           RAM_13_123_port, IN4 => n4582, IN5 => n4458, Q => 
                           n4463);
   U5796 : AO22X1 port map( IN1 => RAM_3_123_port, IN2 => n4615, IN3 => 
                           RAM_2_123_port, IN4 => n4604, Q => n4459);
   U5797 : AO221X1 port map( IN1 => RAM_0_123_port, IN2 => n4637, IN3 => 
                           RAM_1_123_port, IN4 => n4626, IN5 => n4459, Q => 
                           n4462);
   U5798 : AO22X1 port map( IN1 => RAM_7_123_port, IN2 => n4659, IN3 => 
                           RAM_6_123_port, IN4 => n4648, Q => n4460);
   U5799 : AO221X1 port map( IN1 => RAM_4_123_port, IN2 => n4681, IN3 => 
                           RAM_5_123_port, IN4 => n4670, IN5 => n4460, Q => 
                           n4461);
   U5800 : AO22X1 port map( IN1 => RAM_11_124_port, IN2 => n4527, IN3 => 
                           RAM_10_124_port, IN4 => n4516, Q => n4465);
   U5801 : AO221X1 port map( IN1 => RAM_8_124_port, IN2 => n4549, IN3 => 
                           RAM_9_124_port, IN4 => n4538, IN5 => n4465, Q => 
                           n4472);
   U5802 : AO22X1 port map( IN1 => RAM_15_124_port, IN2 => n4571, IN3 => 
                           RAM_14_124_port, IN4 => n4560, Q => n4466);
   U5803 : AO221X1 port map( IN1 => RAM_12_124_port, IN2 => n4593, IN3 => 
                           RAM_13_124_port, IN4 => n4582, IN5 => n4466, Q => 
                           n4471);
   U5804 : AO22X1 port map( IN1 => RAM_3_124_port, IN2 => n4615, IN3 => 
                           RAM_2_124_port, IN4 => n4604, Q => n4467);
   U5805 : AO221X1 port map( IN1 => RAM_0_124_port, IN2 => n4637, IN3 => 
                           RAM_1_124_port, IN4 => n4626, IN5 => n4467, Q => 
                           n4470);
   U5806 : AO22X1 port map( IN1 => RAM_7_124_port, IN2 => n4659, IN3 => 
                           RAM_6_124_port, IN4 => n4648, Q => n4468);
   U5807 : AO221X1 port map( IN1 => RAM_4_124_port, IN2 => n4681, IN3 => 
                           RAM_5_124_port, IN4 => n4670, IN5 => n4468, Q => 
                           n4469);
   U5808 : OR4X1 port map( IN1 => n4472, IN2 => n4471, IN3 => n4470, IN4 => 
                           n4469, Q => RAMDOUT2(124));
   U5809 : AO22X1 port map( IN1 => RAM_11_125_port, IN2 => n4527, IN3 => 
                           RAM_10_125_port, IN4 => n4516, Q => n4473);
   U5810 : AO221X1 port map( IN1 => RAM_8_125_port, IN2 => n4549, IN3 => 
                           RAM_9_125_port, IN4 => n4538, IN5 => n4473, Q => 
                           n4480);
   U5811 : AO22X1 port map( IN1 => RAM_15_125_port, IN2 => n4571, IN3 => 
                           RAM_14_125_port, IN4 => n4560, Q => n4474);
   U5812 : AO221X1 port map( IN1 => RAM_12_125_port, IN2 => n4593, IN3 => 
                           RAM_13_125_port, IN4 => n4582, IN5 => n4474, Q => 
                           n4479);
   U5813 : AO22X1 port map( IN1 => RAM_3_125_port, IN2 => n4615, IN3 => 
                           RAM_2_125_port, IN4 => n4604, Q => n4475);
   U5814 : AO221X1 port map( IN1 => RAM_0_125_port, IN2 => n4637, IN3 => 
                           RAM_1_125_port, IN4 => n4626, IN5 => n4475, Q => 
                           n4478);
   U5815 : AO22X1 port map( IN1 => RAM_7_125_port, IN2 => n4659, IN3 => 
                           RAM_6_125_port, IN4 => n4648, Q => n4476);
   U5816 : AO221X1 port map( IN1 => RAM_4_125_port, IN2 => n4681, IN3 => 
                           RAM_5_125_port, IN4 => n4670, IN5 => n4476, Q => 
                           n4477);
   U5817 : OR4X1 port map( IN1 => n4480, IN2 => n4479, IN3 => n4478, IN4 => 
                           n4477, Q => RAMDOUT2(125));
   U5818 : AO22X1 port map( IN1 => RAM_11_126_port, IN2 => n4527, IN3 => 
                           RAM_10_126_port, IN4 => n4516, Q => n4481);
   U5819 : AO221X1 port map( IN1 => RAM_8_126_port, IN2 => n4549, IN3 => 
                           RAM_9_126_port, IN4 => n4538, IN5 => n4481, Q => 
                           n4488);
   U5820 : AO22X1 port map( IN1 => RAM_15_126_port, IN2 => n4571, IN3 => 
                           RAM_14_126_port, IN4 => n4560, Q => n4482);
   U5821 : AO221X1 port map( IN1 => RAM_12_126_port, IN2 => n4593, IN3 => 
                           RAM_13_126_port, IN4 => n4582, IN5 => n4482, Q => 
                           n4487);
   U5822 : AO22X1 port map( IN1 => RAM_3_126_port, IN2 => n4615, IN3 => 
                           RAM_2_126_port, IN4 => n4604, Q => n4483);
   U5823 : AO221X1 port map( IN1 => RAM_0_126_port, IN2 => n4637, IN3 => 
                           RAM_1_126_port, IN4 => n4626, IN5 => n4483, Q => 
                           n4486);
   U5824 : AO22X1 port map( IN1 => RAM_7_126_port, IN2 => n4659, IN3 => 
                           RAM_6_126_port, IN4 => n4648, Q => n4484);
   U5825 : AO221X1 port map( IN1 => RAM_4_126_port, IN2 => n4681, IN3 => 
                           RAM_5_126_port, IN4 => n4670, IN5 => n4484, Q => 
                           n4485);
   U5826 : OR4X1 port map( IN1 => n4488, IN2 => n4487, IN3 => n4486, IN4 => 
                           n4485, Q => RAMDOUT2(126));
   U5827 : AO22X1 port map( IN1 => RAM_11_127_port, IN2 => n4527, IN3 => 
                           RAM_10_127_port, IN4 => n4516, Q => n4491);
   U5828 : AO221X1 port map( IN1 => RAM_8_127_port, IN2 => n4549, IN3 => 
                           RAM_9_127_port, IN4 => n4538, IN5 => n4491, Q => 
                           n4512);
   U5829 : AO22X1 port map( IN1 => RAM_15_127_port, IN2 => n4571, IN3 => 
                           RAM_14_127_port, IN4 => n4560, Q => n4496);
   U5830 : AO221X1 port map( IN1 => RAM_12_127_port, IN2 => n4593, IN3 => 
                           RAM_13_127_port, IN4 => n4582, IN5 => n4496, Q => 
                           n4511);
   U5831 : AO22X1 port map( IN1 => RAM_3_127_port, IN2 => n4615, IN3 => 
                           RAM_2_127_port, IN4 => n4604, Q => n4501);
   U5832 : AO221X1 port map( IN1 => RAM_0_127_port, IN2 => n4637, IN3 => 
                           RAM_1_127_port, IN4 => n4626, IN5 => n4501, Q => 
                           n4510);
   U5833 : AO22X1 port map( IN1 => RAM_7_127_port, IN2 => n4659, IN3 => 
                           RAM_6_127_port, IN4 => n4648, Q => n4506);
   U5834 : AO221X1 port map( IN1 => RAM_4_127_port, IN2 => n4681, IN3 => 
                           RAM_5_127_port, IN4 => n4670, IN5 => n4506, Q => 
                           n4509);
   U5835 : OR4X1 port map( IN1 => n4512, IN2 => n4511, IN3 => n4510, IN4 => 
                           n4509, Q => RAMDOUT2(127));
   U5836 : AND2X2 port map( IN1 => n3465, IN2 => n3471, Q => n4493);
   U5837 : AND2X2 port map( IN1 => n3465, IN2 => n3472, Q => n4492);
   U5838 : AND2X2 port map( IN1 => n3465, IN2 => n3473, Q => n4490);
   U5839 : AND2X2 port map( IN1 => n3465, IN2 => n3474, Q => n4489);
   U5840 : AND2X2 port map( IN1 => n3471, IN2 => n3467, Q => n4498);
   U5841 : AND2X2 port map( IN1 => n3472, IN2 => n3467, Q => n4497);
   U5842 : AND2X2 port map( IN1 => n3467, IN2 => n3473, Q => n4495);
   U5843 : AND2X2 port map( IN1 => n3474, IN2 => n3467, Q => n4494);
   U5844 : AND2X2 port map( IN1 => n3469, IN2 => n3471, Q => n4503);
   U5845 : AND2X2 port map( IN1 => n3469, IN2 => n3472, Q => n4502);
   U5846 : AND2X2 port map( IN1 => n3469, IN2 => n3473, Q => n4500);
   U5847 : AND2X2 port map( IN1 => n3469, IN2 => n3474, Q => n4499);
   U5848 : AND2X2 port map( IN1 => n3475, IN2 => n3471, Q => n4508);
   U5849 : AND2X2 port map( IN1 => n3475, IN2 => n3472, Q => n4507);
   U5850 : AND2X2 port map( IN1 => n3475, IN2 => n3473, Q => n4505);
   U5851 : AND2X2 port map( IN1 => n3475, IN2 => n3474, Q => n4504);
   U5852 : INVX0 port map( INP => n29, ZN => n5424);
   U5853 : INVX0 port map( INP => n5341, ZN => n5334);
   U5854 : INVX0 port map( INP => n32, ZN => n5341);
   U5855 : NAND2X0 port map( IN1 => n27, IN2 => n23, QN => n26);
   U5856 : NOR2X0 port map( IN1 => n2496, IN2 => n2810, QN => n30);
   U5857 : NOR2X0 port map( IN1 => n2497, IN2 => n2810, QN => n33);
   U5858 : NAND2X0 port map( IN1 => n25, IN2 => n22, QN => n24);
   U5859 : NAND2X0 port map( IN1 => n27, IN2 => n25, QN => n28);
   U5860 : NAND2X0 port map( IN1 => n30, IN2 => n25, QN => n31);
   U5861 : NAND2X0 port map( IN1 => n33, IN2 => n25, QN => n35);
   U5862 : INVX0 port map( INP => n24, ZN => n5548);
   U5863 : AND2X1 port map( IN1 => RAMWRITE1, IN2 => RAMADDR1(3), Q => n34);
   U5864 : NOR2X0 port map( IN1 => n5616, IN2 => n2496, QN => n22);
   U5865 : INVX0 port map( INP => RAMADDR1(0), ZN => n5615);
   U5866 : NAND2X0 port map( IN1 => n37, IN2 => n30, QN => n42);
   U5867 : NAND2X0 port map( IN1 => n37, IN2 => n22, QN => n36);
   U5868 : NAND2X0 port map( IN1 => n37, IN2 => n33, QN => n44);
   U5869 : NAND2X0 port map( IN1 => n37, IN2 => n27, QN => n40);
   U5870 : NAND2X0 port map( IN1 => n39, IN2 => n30, QN => n43);
   U5871 : NAND2X0 port map( IN1 => n39, IN2 => n22, QN => n38);
   U5872 : NAND2X0 port map( IN1 => n39, IN2 => n33, QN => n46);
   U5873 : NAND2X0 port map( IN1 => n39, IN2 => n27, QN => n41);
   U5874 : NOR2X0 port map( IN1 => n5617, IN2 => RAMADDR1(3), QN => n45);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_LWC_1.all;

entity DATA_PISO_1 is

   port( clk, rst : in std_logic;  data_size_p : in std_logic_vector (2 downto 
         0);  data_size_s : out std_logic_vector (2 downto 0);  data_s : out 
         std_logic_vector (31 downto 0);  data_valid_s : out std_logic;  
         data_ready_s : in std_logic;  data_p : in std_logic_vector (31 downto 
         0);  data_valid_p : in std_logic;  data_ready_p : out std_logic;  
         valid_bytes_p : in std_logic_vector (3 downto 0);  valid_bytes_s : out
         std_logic_vector (3 downto 0);  pad_loc_p : in std_logic_vector (3 
         downto 0);  pad_loc_s : out std_logic_vector (3 downto 0);  eoi_p : in
         std_logic;  eoi_s : out std_logic;  eot_p : in std_logic;  eot_s : out
         std_logic);

end DATA_PISO_1;

architecture SYN_behavioral of DATA_PISO_1 is

begin
   data_size_s <= ( data_size_p(2), data_size_p(1), data_size_p(0) );
   data_s <= ( data_p(31), data_p(30), data_p(29), data_p(28), data_p(27), 
      data_p(26), data_p(25), data_p(24), data_p(23), data_p(22), data_p(21), 
      data_p(20), data_p(19), data_p(18), data_p(17), data_p(16), data_p(15), 
      data_p(14), data_p(13), data_p(12), data_p(11), data_p(10), data_p(9), 
      data_p(8), data_p(7), data_p(6), data_p(5), data_p(4), data_p(3), 
      data_p(2), data_p(1), data_p(0) );
   data_valid_s <= data_valid_p;
   data_ready_p <= data_ready_s;
   valid_bytes_s <= ( valid_bytes_p(3), valid_bytes_p(2), valid_bytes_p(1), 
      valid_bytes_p(0) );
   pad_loc_s <= ( pad_loc_p(3), pad_loc_p(2), pad_loc_p(1), pad_loc_p(0) );
   eoi_s <= eoi_p;
   eot_s <= eot_p;

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_LWC_1.all;

entity KEY_PISO_1 is

   port( clk, rst : in std_logic;  data_s : out std_logic_vector (31 downto 0);
         data_valid_s : out std_logic;  data_ready_s : in std_logic;  data_p : 
         in std_logic_vector (31 downto 0);  data_valid_p : in std_logic;  
         data_ready_p : out std_logic);

end KEY_PISO_1;

architecture SYN_behavioral of KEY_PISO_1 is

begin
   data_s <= ( data_p(31), data_p(30), data_p(29), data_p(28), data_p(27), 
      data_p(26), data_p(25), data_p(24), data_p(23), data_p(22), data_p(21), 
      data_p(20), data_p(19), data_p(18), data_p(17), data_p(16), data_p(15), 
      data_p(14), data_p(13), data_p(12), data_p(11), data_p(10), data_p(9), 
      data_p(8), data_p(7), data_p(6), data_p(5), data_p(4), data_p(3), 
      data_p(2), data_p(1), data_p(0) );
   data_valid_s <= data_valid_p;
   data_ready_p <= data_ready_s;

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_LWC_1.all;

entity StepDownCountLd_N16_step4_1_0 is

   port( clk, len, ena : in std_logic;  load : in std_logic_vector (15 downto 
         0);  count : out std_logic_vector (15 downto 0));

end StepDownCountLd_N16_step4_1_0;

architecture SYN_StepDownCountLd of StepDownCountLd_N16_step4_1_0 is

   component XNOR2X1
      port( IN1, IN2 : in std_logic;  Q : out std_logic);
   end component;
   
   component OR2X1
      port( IN1, IN2 : in std_logic;  Q : out std_logic);
   end component;
   
   component NOR2X0
      port( IN1, IN2 : in std_logic;  QN : out std_logic);
   end component;
   
   component NBUFFX2
      port( INP : in std_logic;  Z : out std_logic);
   end component;
   
   component AO222X1
      port( IN1, IN2, IN3, IN4, IN5, IN6 : in std_logic;  Q : out std_logic);
   end component;
   
   component DFFX1
      port( D, CLK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal count_15_port, count_14_port, count_13_port, count_12_port, 
      count_11_port, count_10_port, count_9_port, count_8_port, count_7_port, 
      count_6_port, count_5_port, count_4_port, count_3_port, count_2_port, N4,
      N5, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18, N19, n3, 
      n4_port, n5_port, n6, n7_port, n8_port, n9_port, n10_port, n11_port, 
      n12_port, n13_port, n14_port, n15_port, n16_port, n17_port, n18_port, 
      n19_port, n20, sub_55_carry_4_port, sub_55_carry_5_port, 
      sub_55_carry_6_port, sub_55_carry_7_port, sub_55_carry_8_port, 
      sub_55_carry_9_port, sub_55_carry_10_port, sub_55_carry_11_port, 
      sub_55_carry_12_port, sub_55_carry_13_port, sub_55_carry_14_port, n1, n2,
      n21, n22, n23, n_3077, n_3078, n_3079, n_3080, n_3081, n_3082, n_3083, 
      n_3084, n_3085, n_3086, n_3087, n_3088, n_3089, n_3090 : std_logic;

begin
   count <= ( count_15_port, count_14_port, count_13_port, count_12_port, 
      count_11_port, count_10_port, count_9_port, count_8_port, count_7_port, 
      count_6_port, count_5_port, count_4_port, count_3_port, count_2_port, N5,
      N4 );
   
   qtemp_reg_0_inst : DFFX1 port map( D => n20, CLK => clk, Q => N4, QN => 
                           n_3077);
   qtemp_reg_1_inst : DFFX1 port map( D => n19_port, CLK => clk, Q => N5, QN =>
                           n_3078);
   qtemp_reg_2_inst : DFFX1 port map( D => n18_port, CLK => clk, Q => 
                           count_2_port, QN => n1);
   qtemp_reg_3_inst : DFFX1 port map( D => n17_port, CLK => clk, Q => 
                           count_3_port, QN => n_3079);
   qtemp_reg_4_inst : DFFX1 port map( D => n16_port, CLK => clk, Q => 
                           count_4_port, QN => n_3080);
   qtemp_reg_5_inst : DFFX1 port map( D => n15_port, CLK => clk, Q => 
                           count_5_port, QN => n_3081);
   qtemp_reg_6_inst : DFFX1 port map( D => n14_port, CLK => clk, Q => 
                           count_6_port, QN => n_3082);
   qtemp_reg_7_inst : DFFX1 port map( D => n13_port, CLK => clk, Q => 
                           count_7_port, QN => n_3083);
   qtemp_reg_8_inst : DFFX1 port map( D => n12_port, CLK => clk, Q => 
                           count_8_port, QN => n_3084);
   qtemp_reg_9_inst : DFFX1 port map( D => n11_port, CLK => clk, Q => 
                           count_9_port, QN => n_3085);
   qtemp_reg_10_inst : DFFX1 port map( D => n10_port, CLK => clk, Q => 
                           count_10_port, QN => n_3086);
   qtemp_reg_11_inst : DFFX1 port map( D => n9_port, CLK => clk, Q => 
                           count_11_port, QN => n_3087);
   qtemp_reg_12_inst : DFFX1 port map( D => n8_port, CLK => clk, Q => 
                           count_12_port, QN => n_3088);
   qtemp_reg_13_inst : DFFX1 port map( D => n7_port, CLK => clk, Q => 
                           count_13_port, QN => n_3089);
   qtemp_reg_14_inst : DFFX1 port map( D => n6, CLK => clk, Q => count_14_port,
                           QN => n_3090);
   qtemp_reg_15_inst : DFFX1 port map( D => n5_port, CLK => clk, Q => 
                           count_15_port, QN => n21);
   U6 : AO222X1 port map( IN1 => load(15), IN2 => n23, IN3 => N19, IN4 => n3, 
                           IN5 => count_15_port, IN6 => n4_port, Q => n5_port);
   U7 : AO222X1 port map( IN1 => load(14), IN2 => n23, IN3 => N18, IN4 => n3, 
                           IN5 => count_14_port, IN6 => n4_port, Q => n6);
   U8 : AO222X1 port map( IN1 => load(13), IN2 => n23, IN3 => N17, IN4 => n3, 
                           IN5 => count_13_port, IN6 => n4_port, Q => n7_port);
   U9 : AO222X1 port map( IN1 => load(12), IN2 => n23, IN3 => N16, IN4 => n3, 
                           IN5 => count_12_port, IN6 => n4_port, Q => n8_port);
   U10 : AO222X1 port map( IN1 => load(11), IN2 => n23, IN3 => N15, IN4 => n3, 
                           IN5 => count_11_port, IN6 => n4_port, Q => n9_port);
   U11 : AO222X1 port map( IN1 => load(10), IN2 => n23, IN3 => N14, IN4 => n3, 
                           IN5 => count_10_port, IN6 => n4_port, Q => n10_port)
                           ;
   U12 : AO222X1 port map( IN1 => load(9), IN2 => n23, IN3 => N13, IN4 => n3, 
                           IN5 => count_9_port, IN6 => n4_port, Q => n11_port);
   U13 : AO222X1 port map( IN1 => load(8), IN2 => n23, IN3 => N12, IN4 => n3, 
                           IN5 => count_8_port, IN6 => n4_port, Q => n12_port);
   U14 : AO222X1 port map( IN1 => load(7), IN2 => n23, IN3 => N11, IN4 => n3, 
                           IN5 => count_7_port, IN6 => n4_port, Q => n13_port);
   U15 : AO222X1 port map( IN1 => load(6), IN2 => n23, IN3 => N10, IN4 => n3, 
                           IN5 => count_6_port, IN6 => n4_port, Q => n14_port);
   U16 : AO222X1 port map( IN1 => load(5), IN2 => n23, IN3 => N9, IN4 => n3, 
                           IN5 => count_5_port, IN6 => n4_port, Q => n15_port);
   U17 : AO222X1 port map( IN1 => load(4), IN2 => n23, IN3 => N8, IN4 => n3, 
                           IN5 => count_4_port, IN6 => n4_port, Q => n16_port);
   U18 : AO222X1 port map( IN1 => load(3), IN2 => n23, IN3 => N7, IN4 => n3, 
                           IN5 => count_3_port, IN6 => n4_port, Q => n17_port);
   U19 : AO222X1 port map( IN1 => load(2), IN2 => n23, IN3 => n1, IN4 => n3, 
                           IN5 => count_2_port, IN6 => n4_port, Q => n18_port);
   U20 : AO222X1 port map( IN1 => load(1), IN2 => n23, IN3 => N5, IN4 => n3, 
                           IN5 => N5, IN6 => n4_port, Q => n19_port);
   U21 : AO222X1 port map( IN1 => load(0), IN2 => n23, IN3 => N4, IN4 => n3, 
                           IN5 => N4, IN6 => n4_port, Q => n20);
   U3 : NOR2X0 port map( IN1 => n4_port, IN2 => n22, QN => n3);
   U4 : NBUFFX2 port map( INP => len, Z => n22);
   U5 : NBUFFX2 port map( INP => len, Z => n23);
   U22 : NOR2X0 port map( IN1 => ena, IN2 => n22, QN => n4_port);
   U23 : XNOR2X1 port map( IN1 => n2, IN2 => n21, Q => N19);
   U24 : NOR2X0 port map( IN1 => sub_55_carry_14_port, IN2 => count_14_port, QN
                           => n2);
   U25 : XNOR2X1 port map( IN1 => count_14_port, IN2 => sub_55_carry_14_port, Q
                           => N18);
   U26 : OR2X1 port map( IN1 => sub_55_carry_13_port, IN2 => count_13_port, Q 
                           => sub_55_carry_14_port);
   U27 : XNOR2X1 port map( IN1 => count_13_port, IN2 => sub_55_carry_13_port, Q
                           => N17);
   U28 : OR2X1 port map( IN1 => sub_55_carry_12_port, IN2 => count_12_port, Q 
                           => sub_55_carry_13_port);
   U29 : XNOR2X1 port map( IN1 => count_12_port, IN2 => sub_55_carry_12_port, Q
                           => N16);
   U30 : OR2X1 port map( IN1 => sub_55_carry_11_port, IN2 => count_11_port, Q 
                           => sub_55_carry_12_port);
   U31 : XNOR2X1 port map( IN1 => count_11_port, IN2 => sub_55_carry_11_port, Q
                           => N15);
   U32 : OR2X1 port map( IN1 => sub_55_carry_10_port, IN2 => count_10_port, Q 
                           => sub_55_carry_11_port);
   U33 : XNOR2X1 port map( IN1 => count_10_port, IN2 => sub_55_carry_10_port, Q
                           => N14);
   U34 : OR2X1 port map( IN1 => sub_55_carry_9_port, IN2 => count_9_port, Q => 
                           sub_55_carry_10_port);
   U35 : XNOR2X1 port map( IN1 => count_9_port, IN2 => sub_55_carry_9_port, Q 
                           => N13);
   U36 : OR2X1 port map( IN1 => sub_55_carry_8_port, IN2 => count_8_port, Q => 
                           sub_55_carry_9_port);
   U37 : XNOR2X1 port map( IN1 => count_8_port, IN2 => sub_55_carry_8_port, Q 
                           => N12);
   U38 : OR2X1 port map( IN1 => sub_55_carry_7_port, IN2 => count_7_port, Q => 
                           sub_55_carry_8_port);
   U39 : XNOR2X1 port map( IN1 => count_7_port, IN2 => sub_55_carry_7_port, Q 
                           => N11);
   U40 : OR2X1 port map( IN1 => sub_55_carry_6_port, IN2 => count_6_port, Q => 
                           sub_55_carry_7_port);
   U41 : XNOR2X1 port map( IN1 => count_6_port, IN2 => sub_55_carry_6_port, Q 
                           => N10);
   U42 : OR2X1 port map( IN1 => sub_55_carry_5_port, IN2 => count_5_port, Q => 
                           sub_55_carry_6_port);
   U43 : XNOR2X1 port map( IN1 => count_5_port, IN2 => sub_55_carry_5_port, Q 
                           => N9);
   U44 : OR2X1 port map( IN1 => sub_55_carry_4_port, IN2 => count_4_port, Q => 
                           sub_55_carry_5_port);
   U45 : XNOR2X1 port map( IN1 => count_4_port, IN2 => sub_55_carry_4_port, Q 
                           => N8);
   U46 : OR2X1 port map( IN1 => count_2_port, IN2 => count_3_port, Q => 
                           sub_55_carry_4_port);
   U47 : XNOR2X1 port map( IN1 => count_3_port, IN2 => count_2_port, Q => N7);

end SYN_StepDownCountLd;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_LWC_1.all;

entity fwft_fifo_G_W32_G_LOG2DEPTH2 is

   port( clk, rst : in std_logic;  din : in std_logic_vector (31 downto 0);  
         din_valid : in std_logic;  din_ready : out std_logic;  dout : out 
         std_logic_vector (31 downto 0);  dout_valid : out std_logic;  
         dout_ready : in std_logic);

end fwft_fifo_G_W32_G_LOG2DEPTH2;

architecture SYN_structure of fwft_fifo_G_W32_G_LOG2DEPTH2 is

   component AO221X1
      port( IN1, IN2, IN3, IN4, IN5 : in std_logic;  Q : out std_logic);
   end component;
   
   component AO22X1
      port( IN1, IN2, IN3, IN4 : in std_logic;  Q : out std_logic);
   end component;
   
   component NOR2X0
      port( IN1, IN2 : in std_logic;  QN : out std_logic);
   end component;
   
   component NBUFFX2
      port( INP : in std_logic;  Z : out std_logic);
   end component;
   
   component INVX0
      port( INP : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2X1
      port( IN1, IN2 : in std_logic;  QN : out std_logic);
   end component;
   
   component NAND3X0
      port( IN1, IN2, IN3 : in std_logic;  QN : out std_logic);
   end component;
   
   component AO21X1
      port( IN1, IN2, IN3 : in std_logic;  Q : out std_logic);
   end component;
   
   component XOR2X1
      port( IN1, IN2 : in std_logic;  Q : out std_logic);
   end component;
   
   component OA21X1
      port( IN1, IN2, IN3 : in std_logic;  Q : out std_logic);
   end component;
   
   component OAI22X1
      port( IN1, IN2, IN3, IN4 : in std_logic;  QN : out std_logic);
   end component;
   
   component AND3X1
      port( IN1, IN2, IN3 : in std_logic;  Q : out std_logic);
   end component;
   
   component OR2X1
      port( IN1, IN2 : in std_logic;  Q : out std_logic);
   end component;
   
   component NAND4X0
      port( IN1, IN2, IN3, IN4 : in std_logic;  QN : out std_logic);
   end component;
   
   component DFFX1
      port( D, CLK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal N10, N11, mem_s_0_31_port, mem_s_0_30_port, mem_s_0_29_port, 
      mem_s_0_28_port, mem_s_0_27_port, mem_s_0_26_port, mem_s_0_25_port, 
      mem_s_0_24_port, mem_s_0_23_port, mem_s_0_22_port, mem_s_0_21_port, 
      mem_s_0_20_port, mem_s_0_19_port, mem_s_0_18_port, mem_s_0_17_port, 
      mem_s_0_16_port, mem_s_0_15_port, mem_s_0_14_port, mem_s_0_13_port, 
      mem_s_0_12_port, mem_s_0_11_port, mem_s_0_10_port, mem_s_0_9_port, 
      mem_s_0_8_port, mem_s_0_7_port, mem_s_0_6_port, mem_s_0_5_port, 
      mem_s_0_4_port, mem_s_0_3_port, mem_s_0_2_port, mem_s_0_1_port, 
      mem_s_0_0_port, mem_s_1_31_port, mem_s_1_30_port, mem_s_1_29_port, 
      mem_s_1_28_port, mem_s_1_27_port, mem_s_1_26_port, mem_s_1_25_port, 
      mem_s_1_24_port, mem_s_1_23_port, mem_s_1_22_port, mem_s_1_21_port, 
      mem_s_1_20_port, mem_s_1_19_port, mem_s_1_18_port, mem_s_1_17_port, 
      mem_s_1_16_port, mem_s_1_15_port, mem_s_1_14_port, mem_s_1_13_port, 
      mem_s_1_12_port, mem_s_1_11_port, mem_s_1_10_port, mem_s_1_9_port, 
      mem_s_1_8_port, mem_s_1_7_port, mem_s_1_6_port, mem_s_1_5_port, 
      mem_s_1_4_port, mem_s_1_3_port, mem_s_1_2_port, mem_s_1_1_port, 
      mem_s_1_0_port, mem_s_2_31_port, mem_s_2_30_port, mem_s_2_29_port, 
      mem_s_2_28_port, mem_s_2_27_port, mem_s_2_26_port, mem_s_2_25_port, 
      mem_s_2_24_port, mem_s_2_23_port, mem_s_2_22_port, mem_s_2_21_port, 
      mem_s_2_20_port, mem_s_2_19_port, mem_s_2_18_port, mem_s_2_17_port, 
      mem_s_2_16_port, mem_s_2_15_port, mem_s_2_14_port, mem_s_2_13_port, 
      mem_s_2_12_port, mem_s_2_11_port, mem_s_2_10_port, mem_s_2_9_port, 
      mem_s_2_8_port, mem_s_2_7_port, mem_s_2_6_port, mem_s_2_5_port, 
      mem_s_2_4_port, mem_s_2_3_port, mem_s_2_2_port, mem_s_2_1_port, 
      mem_s_2_0_port, mem_s_3_31_port, mem_s_3_30_port, mem_s_3_29_port, 
      mem_s_3_28_port, mem_s_3_27_port, mem_s_3_26_port, mem_s_3_25_port, 
      mem_s_3_24_port, mem_s_3_23_port, mem_s_3_22_port, mem_s_3_21_port, 
      mem_s_3_20_port, mem_s_3_19_port, mem_s_3_18_port, mem_s_3_17_port, 
      mem_s_3_16_port, mem_s_3_15_port, mem_s_3_14_port, mem_s_3_13_port, 
      mem_s_3_12_port, mem_s_3_11_port, mem_s_3_10_port, mem_s_3_9_port, 
      mem_s_3_8_port, mem_s_3_7_port, mem_s_3_6_port, mem_s_3_5_port, 
      mem_s_3_4_port, mem_s_3_3_port, mem_s_3_2_port, mem_s_3_1_port, 
      mem_s_3_0_port, entries_s_1_port, entries_s_0_port, N12, wr_ptr_s_1_port,
      wr_ptr_s_0_port, n13, n14, din_ready_port, n21, n22, n24, n25, n26, n27, 
      n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42
      , n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, 
      n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71
      , n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, 
      n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, 
      n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, 
      n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, 
      n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, 
      n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, 
      n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, 
      n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, 
      n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, 
      dout_valid_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10_port, n11_port, 
      n12_port, n15, n16, n17, n18, n19, n20, n23, n184, n185, n186, n187, n188
      , n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
      n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, 
      n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, 
      n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, 
      n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, 
      n249, n250, n251, n_3091, n_3092, n_3093, n_3094, n_3095, n_3096, n_3097,
      n_3098, n_3099, n_3100, n_3101, n_3102, n_3103, n_3104, n_3105, n_3106, 
      n_3107, n_3108, n_3109, n_3110, n_3111, n_3112, n_3113, n_3114, n_3115, 
      n_3116, n_3117, n_3118, n_3119, n_3120, n_3121, n_3122, n_3123, n_3124, 
      n_3125, n_3126, n_3127, n_3128, n_3129, n_3130, n_3131, n_3132, n_3133, 
      n_3134, n_3135, n_3136, n_3137, n_3138, n_3139, n_3140, n_3141, n_3142, 
      n_3143, n_3144, n_3145, n_3146, n_3147, n_3148, n_3149, n_3150, n_3151, 
      n_3152, n_3153, n_3154, n_3155, n_3156, n_3157, n_3158, n_3159, n_3160, 
      n_3161, n_3162, n_3163, n_3164, n_3165, n_3166, n_3167, n_3168, n_3169, 
      n_3170, n_3171, n_3172, n_3173, n_3174, n_3175, n_3176, n_3177, n_3178, 
      n_3179, n_3180, n_3181, n_3182, n_3183, n_3184, n_3185, n_3186, n_3187, 
      n_3188, n_3189, n_3190, n_3191, n_3192, n_3193, n_3194, n_3195, n_3196, 
      n_3197, n_3198, n_3199, n_3200, n_3201, n_3202, n_3203, n_3204, n_3205, 
      n_3206, n_3207, n_3208, n_3209, n_3210, n_3211, n_3212, n_3213, n_3214, 
      n_3215, n_3216, n_3217, n_3218, n_3219 : std_logic;

begin
   din_ready <= din_ready_port;
   dout_valid <= dout_valid_port;
   
   entries_s_reg_0_inst : DFFX1 port map( D => n183, CLK => n214, Q => 
                           entries_s_0_port, QN => n22);
   entries_s_reg_2_inst : DFFX1 port map( D => n179, CLK => n214, Q => N12, QN 
                           => din_ready_port);
   entries_s_reg_1_inst : DFFX1 port map( D => n180, CLK => n214, Q => 
                           entries_s_1_port, QN => n21);
   rd_ptr_s_reg_0_inst : DFFX1 port map( D => n181, CLK => n214, Q => N10, QN 
                           => n14);
   rd_ptr_s_reg_1_inst : DFFX1 port map( D => n182, CLK => n214, Q => N11, QN 
                           => n1);
   wr_ptr_s_reg_0_inst : DFFX1 port map( D => n177, CLK => n214, Q => 
                           wr_ptr_s_0_port, QN => n_3091);
   wr_ptr_s_reg_1_inst : DFFX1 port map( D => n178, CLK => n214, Q => 
                           wr_ptr_s_1_port, QN => n13);
   mem_s_reg_3_0_inst : DFFX1 port map( D => n176, CLK => n214, Q => 
                           mem_s_3_0_port, QN => n_3092);
   mem_s_reg_3_1_inst : DFFX1 port map( D => n175, CLK => n214, Q => 
                           mem_s_3_1_port, QN => n_3093);
   mem_s_reg_3_2_inst : DFFX1 port map( D => n174, CLK => n214, Q => 
                           mem_s_3_2_port, QN => n_3094);
   mem_s_reg_3_3_inst : DFFX1 port map( D => n173, CLK => n214, Q => 
                           mem_s_3_3_port, QN => n_3095);
   mem_s_reg_3_4_inst : DFFX1 port map( D => n172, CLK => n214, Q => 
                           mem_s_3_4_port, QN => n_3096);
   mem_s_reg_3_5_inst : DFFX1 port map( D => n171, CLK => n215, Q => 
                           mem_s_3_5_port, QN => n_3097);
   mem_s_reg_3_6_inst : DFFX1 port map( D => n170, CLK => n215, Q => 
                           mem_s_3_6_port, QN => n_3098);
   mem_s_reg_3_7_inst : DFFX1 port map( D => n169, CLK => n215, Q => 
                           mem_s_3_7_port, QN => n_3099);
   mem_s_reg_3_8_inst : DFFX1 port map( D => n168, CLK => n215, Q => 
                           mem_s_3_8_port, QN => n_3100);
   mem_s_reg_3_9_inst : DFFX1 port map( D => n167, CLK => n215, Q => 
                           mem_s_3_9_port, QN => n_3101);
   mem_s_reg_3_10_inst : DFFX1 port map( D => n166, CLK => n215, Q => 
                           mem_s_3_10_port, QN => n_3102);
   mem_s_reg_3_11_inst : DFFX1 port map( D => n165, CLK => n215, Q => 
                           mem_s_3_11_port, QN => n_3103);
   mem_s_reg_3_12_inst : DFFX1 port map( D => n164, CLK => n215, Q => 
                           mem_s_3_12_port, QN => n_3104);
   mem_s_reg_3_13_inst : DFFX1 port map( D => n163, CLK => n215, Q => 
                           mem_s_3_13_port, QN => n_3105);
   mem_s_reg_3_14_inst : DFFX1 port map( D => n162, CLK => n215, Q => 
                           mem_s_3_14_port, QN => n_3106);
   mem_s_reg_3_15_inst : DFFX1 port map( D => n161, CLK => n215, Q => 
                           mem_s_3_15_port, QN => n_3107);
   mem_s_reg_3_16_inst : DFFX1 port map( D => n160, CLK => n215, Q => 
                           mem_s_3_16_port, QN => n_3108);
   mem_s_reg_3_17_inst : DFFX1 port map( D => n159, CLK => n216, Q => 
                           mem_s_3_17_port, QN => n_3109);
   mem_s_reg_3_18_inst : DFFX1 port map( D => n158, CLK => n216, Q => 
                           mem_s_3_18_port, QN => n_3110);
   mem_s_reg_3_19_inst : DFFX1 port map( D => n157, CLK => n216, Q => 
                           mem_s_3_19_port, QN => n_3111);
   mem_s_reg_3_20_inst : DFFX1 port map( D => n156, CLK => n216, Q => 
                           mem_s_3_20_port, QN => n_3112);
   mem_s_reg_3_21_inst : DFFX1 port map( D => n155, CLK => n216, Q => 
                           mem_s_3_21_port, QN => n_3113);
   mem_s_reg_3_22_inst : DFFX1 port map( D => n154, CLK => n216, Q => 
                           mem_s_3_22_port, QN => n_3114);
   mem_s_reg_3_23_inst : DFFX1 port map( D => n153, CLK => n216, Q => 
                           mem_s_3_23_port, QN => n_3115);
   mem_s_reg_3_24_inst : DFFX1 port map( D => n152, CLK => n216, Q => 
                           mem_s_3_24_port, QN => n_3116);
   mem_s_reg_3_25_inst : DFFX1 port map( D => n151, CLK => n216, Q => 
                           mem_s_3_25_port, QN => n_3117);
   mem_s_reg_3_26_inst : DFFX1 port map( D => n150, CLK => n216, Q => 
                           mem_s_3_26_port, QN => n_3118);
   mem_s_reg_3_27_inst : DFFX1 port map( D => n149, CLK => n216, Q => 
                           mem_s_3_27_port, QN => n_3119);
   mem_s_reg_3_28_inst : DFFX1 port map( D => n148, CLK => n216, Q => 
                           mem_s_3_28_port, QN => n_3120);
   mem_s_reg_3_29_inst : DFFX1 port map( D => n147, CLK => n217, Q => 
                           mem_s_3_29_port, QN => n_3121);
   mem_s_reg_3_30_inst : DFFX1 port map( D => n146, CLK => n217, Q => 
                           mem_s_3_30_port, QN => n_3122);
   mem_s_reg_3_31_inst : DFFX1 port map( D => n145, CLK => n217, Q => 
                           mem_s_3_31_port, QN => n_3123);
   mem_s_reg_2_0_inst : DFFX1 port map( D => n144, CLK => n217, Q => 
                           mem_s_2_0_port, QN => n_3124);
   mem_s_reg_2_1_inst : DFFX1 port map( D => n143, CLK => n217, Q => 
                           mem_s_2_1_port, QN => n_3125);
   mem_s_reg_2_2_inst : DFFX1 port map( D => n142, CLK => n217, Q => 
                           mem_s_2_2_port, QN => n_3126);
   mem_s_reg_2_3_inst : DFFX1 port map( D => n141, CLK => n217, Q => 
                           mem_s_2_3_port, QN => n_3127);
   mem_s_reg_2_4_inst : DFFX1 port map( D => n140, CLK => n217, Q => 
                           mem_s_2_4_port, QN => n_3128);
   mem_s_reg_2_5_inst : DFFX1 port map( D => n139, CLK => n217, Q => 
                           mem_s_2_5_port, QN => n_3129);
   mem_s_reg_2_6_inst : DFFX1 port map( D => n138, CLK => n217, Q => 
                           mem_s_2_6_port, QN => n_3130);
   mem_s_reg_2_7_inst : DFFX1 port map( D => n137, CLK => n217, Q => 
                           mem_s_2_7_port, QN => n_3131);
   mem_s_reg_2_8_inst : DFFX1 port map( D => n136, CLK => n217, Q => 
                           mem_s_2_8_port, QN => n_3132);
   mem_s_reg_2_9_inst : DFFX1 port map( D => n135, CLK => n218, Q => 
                           mem_s_2_9_port, QN => n_3133);
   mem_s_reg_2_10_inst : DFFX1 port map( D => n134, CLK => n218, Q => 
                           mem_s_2_10_port, QN => n_3134);
   mem_s_reg_2_11_inst : DFFX1 port map( D => n133, CLK => n218, Q => 
                           mem_s_2_11_port, QN => n_3135);
   mem_s_reg_2_12_inst : DFFX1 port map( D => n132, CLK => n218, Q => 
                           mem_s_2_12_port, QN => n_3136);
   mem_s_reg_2_13_inst : DFFX1 port map( D => n131, CLK => n218, Q => 
                           mem_s_2_13_port, QN => n_3137);
   mem_s_reg_2_14_inst : DFFX1 port map( D => n130, CLK => n218, Q => 
                           mem_s_2_14_port, QN => n_3138);
   mem_s_reg_2_15_inst : DFFX1 port map( D => n129, CLK => n218, Q => 
                           mem_s_2_15_port, QN => n_3139);
   mem_s_reg_2_16_inst : DFFX1 port map( D => n128, CLK => n218, Q => 
                           mem_s_2_16_port, QN => n_3140);
   mem_s_reg_2_17_inst : DFFX1 port map( D => n127, CLK => n218, Q => 
                           mem_s_2_17_port, QN => n_3141);
   mem_s_reg_2_18_inst : DFFX1 port map( D => n126, CLK => n218, Q => 
                           mem_s_2_18_port, QN => n_3142);
   mem_s_reg_2_19_inst : DFFX1 port map( D => n125, CLK => n218, Q => 
                           mem_s_2_19_port, QN => n_3143);
   mem_s_reg_2_20_inst : DFFX1 port map( D => n124, CLK => n218, Q => 
                           mem_s_2_20_port, QN => n_3144);
   mem_s_reg_2_21_inst : DFFX1 port map( D => n123, CLK => n219, Q => 
                           mem_s_2_21_port, QN => n_3145);
   mem_s_reg_2_22_inst : DFFX1 port map( D => n122, CLK => n219, Q => 
                           mem_s_2_22_port, QN => n_3146);
   mem_s_reg_2_23_inst : DFFX1 port map( D => n121, CLK => n219, Q => 
                           mem_s_2_23_port, QN => n_3147);
   mem_s_reg_2_24_inst : DFFX1 port map( D => n120, CLK => n219, Q => 
                           mem_s_2_24_port, QN => n_3148);
   mem_s_reg_2_25_inst : DFFX1 port map( D => n119, CLK => n219, Q => 
                           mem_s_2_25_port, QN => n_3149);
   mem_s_reg_2_26_inst : DFFX1 port map( D => n118, CLK => n219, Q => 
                           mem_s_2_26_port, QN => n_3150);
   mem_s_reg_2_27_inst : DFFX1 port map( D => n117, CLK => n219, Q => 
                           mem_s_2_27_port, QN => n_3151);
   mem_s_reg_2_28_inst : DFFX1 port map( D => n116, CLK => n219, Q => 
                           mem_s_2_28_port, QN => n_3152);
   mem_s_reg_2_29_inst : DFFX1 port map( D => n115, CLK => n219, Q => 
                           mem_s_2_29_port, QN => n_3153);
   mem_s_reg_2_30_inst : DFFX1 port map( D => n114, CLK => n219, Q => 
                           mem_s_2_30_port, QN => n_3154);
   mem_s_reg_2_31_inst : DFFX1 port map( D => n113, CLK => n219, Q => 
                           mem_s_2_31_port, QN => n_3155);
   mem_s_reg_1_0_inst : DFFX1 port map( D => n112, CLK => n219, Q => 
                           mem_s_1_0_port, QN => n_3156);
   mem_s_reg_1_1_inst : DFFX1 port map( D => n111, CLK => n220, Q => 
                           mem_s_1_1_port, QN => n_3157);
   mem_s_reg_1_2_inst : DFFX1 port map( D => n110, CLK => n220, Q => 
                           mem_s_1_2_port, QN => n_3158);
   mem_s_reg_1_3_inst : DFFX1 port map( D => n109, CLK => n220, Q => 
                           mem_s_1_3_port, QN => n_3159);
   mem_s_reg_1_4_inst : DFFX1 port map( D => n108, CLK => n220, Q => 
                           mem_s_1_4_port, QN => n_3160);
   mem_s_reg_1_5_inst : DFFX1 port map( D => n107, CLK => n220, Q => 
                           mem_s_1_5_port, QN => n_3161);
   mem_s_reg_1_6_inst : DFFX1 port map( D => n106, CLK => n220, Q => 
                           mem_s_1_6_port, QN => n_3162);
   mem_s_reg_1_7_inst : DFFX1 port map( D => n105, CLK => n220, Q => 
                           mem_s_1_7_port, QN => n_3163);
   mem_s_reg_1_8_inst : DFFX1 port map( D => n104, CLK => n220, Q => 
                           mem_s_1_8_port, QN => n_3164);
   mem_s_reg_1_9_inst : DFFX1 port map( D => n103, CLK => n220, Q => 
                           mem_s_1_9_port, QN => n_3165);
   mem_s_reg_1_10_inst : DFFX1 port map( D => n102, CLK => n220, Q => 
                           mem_s_1_10_port, QN => n_3166);
   mem_s_reg_1_11_inst : DFFX1 port map( D => n101, CLK => n220, Q => 
                           mem_s_1_11_port, QN => n_3167);
   mem_s_reg_1_12_inst : DFFX1 port map( D => n100, CLK => n220, Q => 
                           mem_s_1_12_port, QN => n_3168);
   mem_s_reg_1_13_inst : DFFX1 port map( D => n99, CLK => n221, Q => 
                           mem_s_1_13_port, QN => n_3169);
   mem_s_reg_1_14_inst : DFFX1 port map( D => n98, CLK => n221, Q => 
                           mem_s_1_14_port, QN => n_3170);
   mem_s_reg_1_15_inst : DFFX1 port map( D => n97, CLK => n221, Q => 
                           mem_s_1_15_port, QN => n_3171);
   mem_s_reg_1_16_inst : DFFX1 port map( D => n96, CLK => n221, Q => 
                           mem_s_1_16_port, QN => n_3172);
   mem_s_reg_1_17_inst : DFFX1 port map( D => n95, CLK => n221, Q => 
                           mem_s_1_17_port, QN => n_3173);
   mem_s_reg_1_18_inst : DFFX1 port map( D => n94, CLK => n221, Q => 
                           mem_s_1_18_port, QN => n_3174);
   mem_s_reg_1_19_inst : DFFX1 port map( D => n93, CLK => n221, Q => 
                           mem_s_1_19_port, QN => n_3175);
   mem_s_reg_1_20_inst : DFFX1 port map( D => n92, CLK => n221, Q => 
                           mem_s_1_20_port, QN => n_3176);
   mem_s_reg_1_21_inst : DFFX1 port map( D => n91, CLK => n221, Q => 
                           mem_s_1_21_port, QN => n_3177);
   mem_s_reg_1_22_inst : DFFX1 port map( D => n90, CLK => n221, Q => 
                           mem_s_1_22_port, QN => n_3178);
   mem_s_reg_1_23_inst : DFFX1 port map( D => n89, CLK => n221, Q => 
                           mem_s_1_23_port, QN => n_3179);
   mem_s_reg_1_24_inst : DFFX1 port map( D => n88, CLK => n221, Q => 
                           mem_s_1_24_port, QN => n_3180);
   mem_s_reg_1_25_inst : DFFX1 port map( D => n87, CLK => n222, Q => 
                           mem_s_1_25_port, QN => n_3181);
   mem_s_reg_1_26_inst : DFFX1 port map( D => n86, CLK => n222, Q => 
                           mem_s_1_26_port, QN => n_3182);
   mem_s_reg_1_27_inst : DFFX1 port map( D => n85, CLK => n222, Q => 
                           mem_s_1_27_port, QN => n_3183);
   mem_s_reg_1_28_inst : DFFX1 port map( D => n84, CLK => n222, Q => 
                           mem_s_1_28_port, QN => n_3184);
   mem_s_reg_1_29_inst : DFFX1 port map( D => n83, CLK => n222, Q => 
                           mem_s_1_29_port, QN => n_3185);
   mem_s_reg_1_30_inst : DFFX1 port map( D => n82, CLK => n222, Q => 
                           mem_s_1_30_port, QN => n_3186);
   mem_s_reg_1_31_inst : DFFX1 port map( D => n81, CLK => n222, Q => 
                           mem_s_1_31_port, QN => n_3187);
   mem_s_reg_0_0_inst : DFFX1 port map( D => n80, CLK => n222, Q => 
                           mem_s_0_0_port, QN => n_3188);
   mem_s_reg_0_1_inst : DFFX1 port map( D => n79, CLK => n222, Q => 
                           mem_s_0_1_port, QN => n_3189);
   mem_s_reg_0_2_inst : DFFX1 port map( D => n78, CLK => n222, Q => 
                           mem_s_0_2_port, QN => n_3190);
   mem_s_reg_0_3_inst : DFFX1 port map( D => n77, CLK => n222, Q => 
                           mem_s_0_3_port, QN => n_3191);
   mem_s_reg_0_4_inst : DFFX1 port map( D => n76, CLK => n222, Q => 
                           mem_s_0_4_port, QN => n_3192);
   mem_s_reg_0_5_inst : DFFX1 port map( D => n75, CLK => n223, Q => 
                           mem_s_0_5_port, QN => n_3193);
   mem_s_reg_0_6_inst : DFFX1 port map( D => n74, CLK => n223, Q => 
                           mem_s_0_6_port, QN => n_3194);
   mem_s_reg_0_7_inst : DFFX1 port map( D => n73, CLK => n223, Q => 
                           mem_s_0_7_port, QN => n_3195);
   mem_s_reg_0_8_inst : DFFX1 port map( D => n72, CLK => n223, Q => 
                           mem_s_0_8_port, QN => n_3196);
   mem_s_reg_0_9_inst : DFFX1 port map( D => n71, CLK => n223, Q => 
                           mem_s_0_9_port, QN => n_3197);
   mem_s_reg_0_10_inst : DFFX1 port map( D => n70, CLK => n223, Q => 
                           mem_s_0_10_port, QN => n_3198);
   mem_s_reg_0_11_inst : DFFX1 port map( D => n69, CLK => n223, Q => 
                           mem_s_0_11_port, QN => n_3199);
   mem_s_reg_0_12_inst : DFFX1 port map( D => n68, CLK => n223, Q => 
                           mem_s_0_12_port, QN => n_3200);
   mem_s_reg_0_13_inst : DFFX1 port map( D => n67, CLK => n223, Q => 
                           mem_s_0_13_port, QN => n_3201);
   mem_s_reg_0_14_inst : DFFX1 port map( D => n66, CLK => n223, Q => 
                           mem_s_0_14_port, QN => n_3202);
   mem_s_reg_0_15_inst : DFFX1 port map( D => n65, CLK => n223, Q => 
                           mem_s_0_15_port, QN => n_3203);
   mem_s_reg_0_16_inst : DFFX1 port map( D => n64, CLK => n223, Q => 
                           mem_s_0_16_port, QN => n_3204);
   mem_s_reg_0_17_inst : DFFX1 port map( D => n63, CLK => n224, Q => 
                           mem_s_0_17_port, QN => n_3205);
   mem_s_reg_0_18_inst : DFFX1 port map( D => n62, CLK => n224, Q => 
                           mem_s_0_18_port, QN => n_3206);
   mem_s_reg_0_19_inst : DFFX1 port map( D => n61, CLK => n224, Q => 
                           mem_s_0_19_port, QN => n_3207);
   mem_s_reg_0_20_inst : DFFX1 port map( D => n60, CLK => n224, Q => 
                           mem_s_0_20_port, QN => n_3208);
   mem_s_reg_0_21_inst : DFFX1 port map( D => n59, CLK => n224, Q => 
                           mem_s_0_21_port, QN => n_3209);
   mem_s_reg_0_22_inst : DFFX1 port map( D => n58, CLK => n224, Q => 
                           mem_s_0_22_port, QN => n_3210);
   mem_s_reg_0_23_inst : DFFX1 port map( D => n57, CLK => n224, Q => 
                           mem_s_0_23_port, QN => n_3211);
   mem_s_reg_0_24_inst : DFFX1 port map( D => n56, CLK => n224, Q => 
                           mem_s_0_24_port, QN => n_3212);
   mem_s_reg_0_25_inst : DFFX1 port map( D => n55, CLK => n224, Q => 
                           mem_s_0_25_port, QN => n_3213);
   mem_s_reg_0_26_inst : DFFX1 port map( D => n54, CLK => n224, Q => 
                           mem_s_0_26_port, QN => n_3214);
   mem_s_reg_0_27_inst : DFFX1 port map( D => n53, CLK => n224, Q => 
                           mem_s_0_27_port, QN => n_3215);
   mem_s_reg_0_28_inst : DFFX1 port map( D => n52, CLK => n224, Q => 
                           mem_s_0_28_port, QN => n_3216);
   mem_s_reg_0_29_inst : DFFX1 port map( D => n51, CLK => n225, Q => 
                           mem_s_0_29_port, QN => n_3217);
   mem_s_reg_0_30_inst : DFFX1 port map( D => n50, CLK => n225, Q => 
                           mem_s_0_30_port, QN => n_3218);
   mem_s_reg_0_31_inst : DFFX1 port map( D => n49, CLK => n225, Q => 
                           mem_s_0_31_port, QN => n_3219);
   U22 : AO22X1 port map( IN1 => din(31), IN2 => n244, IN3 => mem_s_0_31_port, 
                           IN4 => n243, Q => n49);
   U23 : AO22X1 port map( IN1 => din(30), IN2 => n244, IN3 => mem_s_0_30_port, 
                           IN4 => n243, Q => n50);
   U24 : AO22X1 port map( IN1 => din(29), IN2 => n245, IN3 => mem_s_0_29_port, 
                           IN4 => n243, Q => n51);
   U25 : AO22X1 port map( IN1 => din(28), IN2 => n245, IN3 => mem_s_0_28_port, 
                           IN4 => n243, Q => n52);
   U26 : AO22X1 port map( IN1 => din(27), IN2 => n244, IN3 => mem_s_0_27_port, 
                           IN4 => n243, Q => n53);
   U27 : AO22X1 port map( IN1 => din(26), IN2 => n244, IN3 => mem_s_0_26_port, 
                           IN4 => n243, Q => n54);
   U28 : AO22X1 port map( IN1 => din(25), IN2 => n244, IN3 => mem_s_0_25_port, 
                           IN4 => n243, Q => n55);
   U29 : AO22X1 port map( IN1 => din(24), IN2 => n244, IN3 => mem_s_0_24_port, 
                           IN4 => n243, Q => n56);
   U30 : AO22X1 port map( IN1 => din(23), IN2 => n245, IN3 => mem_s_0_23_port, 
                           IN4 => n242, Q => n57);
   U31 : AO22X1 port map( IN1 => din(22), IN2 => n245, IN3 => mem_s_0_22_port, 
                           IN4 => n242, Q => n58);
   U32 : AO22X1 port map( IN1 => din(21), IN2 => n244, IN3 => mem_s_0_21_port, 
                           IN4 => n242, Q => n59);
   U33 : AO22X1 port map( IN1 => din(20), IN2 => n244, IN3 => mem_s_0_20_port, 
                           IN4 => n242, Q => n60);
   U34 : AO22X1 port map( IN1 => din(19), IN2 => n245, IN3 => mem_s_0_19_port, 
                           IN4 => n242, Q => n61);
   U35 : AO22X1 port map( IN1 => din(18), IN2 => n244, IN3 => mem_s_0_18_port, 
                           IN4 => n242, Q => n62);
   U36 : AO22X1 port map( IN1 => din(17), IN2 => n245, IN3 => mem_s_0_17_port, 
                           IN4 => n242, Q => n63);
   U37 : AO22X1 port map( IN1 => din(16), IN2 => n245, IN3 => mem_s_0_16_port, 
                           IN4 => n242, Q => n64);
   U38 : AO22X1 port map( IN1 => din(15), IN2 => n244, IN3 => mem_s_0_15_port, 
                           IN4 => n242, Q => n65);
   U39 : AO22X1 port map( IN1 => din(14), IN2 => n245, IN3 => mem_s_0_14_port, 
                           IN4 => n242, Q => n66);
   U40 : AO22X1 port map( IN1 => din(13), IN2 => n244, IN3 => mem_s_0_13_port, 
                           IN4 => n242, Q => n67);
   U41 : AO22X1 port map( IN1 => din(12), IN2 => n245, IN3 => mem_s_0_12_port, 
                           IN4 => n242, Q => n68);
   U42 : AO22X1 port map( IN1 => din(11), IN2 => n244, IN3 => mem_s_0_11_port, 
                           IN4 => n241, Q => n69);
   U43 : AO22X1 port map( IN1 => din(10), IN2 => n245, IN3 => mem_s_0_10_port, 
                           IN4 => n241, Q => n70);
   U44 : AO22X1 port map( IN1 => din(9), IN2 => n244, IN3 => mem_s_0_9_port, 
                           IN4 => n241, Q => n71);
   U45 : AO22X1 port map( IN1 => din(8), IN2 => n244, IN3 => mem_s_0_8_port, 
                           IN4 => n241, Q => n72);
   U46 : AO22X1 port map( IN1 => din(7), IN2 => n244, IN3 => mem_s_0_7_port, 
                           IN4 => n241, Q => n73);
   U47 : AO22X1 port map( IN1 => din(6), IN2 => n244, IN3 => mem_s_0_6_port, 
                           IN4 => n241, Q => n74);
   U48 : AO22X1 port map( IN1 => din(5), IN2 => n244, IN3 => mem_s_0_5_port, 
                           IN4 => n241, Q => n75);
   U49 : AO22X1 port map( IN1 => din(4), IN2 => n245, IN3 => mem_s_0_4_port, 
                           IN4 => n241, Q => n76);
   U50 : AO22X1 port map( IN1 => din(3), IN2 => n245, IN3 => mem_s_0_3_port, 
                           IN4 => n241, Q => n77);
   U51 : AO22X1 port map( IN1 => din(2), IN2 => n245, IN3 => mem_s_0_2_port, 
                           IN4 => n241, Q => n78);
   U52 : AO22X1 port map( IN1 => din(1), IN2 => n245, IN3 => mem_s_0_1_port, 
                           IN4 => n241, Q => n79);
   U53 : AO22X1 port map( IN1 => din(0), IN2 => n245, IN3 => mem_s_0_0_port, 
                           IN4 => n241, Q => n80);
   U54 : NAND3X0 port map( IN1 => n25, IN2 => n13, IN3 => n249, QN => n24);
   U55 : AO22X1 port map( IN1 => n240, IN2 => din(31), IN3 => mem_s_1_31_port, 
                           IN4 => n238, Q => n81);
   U56 : AO22X1 port map( IN1 => n240, IN2 => din(30), IN3 => mem_s_1_30_port, 
                           IN4 => n238, Q => n82);
   U57 : AO22X1 port map( IN1 => n240, IN2 => din(29), IN3 => mem_s_1_29_port, 
                           IN4 => n238, Q => n83);
   U58 : AO22X1 port map( IN1 => n240, IN2 => din(28), IN3 => mem_s_1_28_port, 
                           IN4 => n238, Q => n84);
   U59 : AO22X1 port map( IN1 => n239, IN2 => din(27), IN3 => mem_s_1_27_port, 
                           IN4 => n238, Q => n85);
   U60 : AO22X1 port map( IN1 => n239, IN2 => din(26), IN3 => mem_s_1_26_port, 
                           IN4 => n238, Q => n86);
   U61 : AO22X1 port map( IN1 => n239, IN2 => din(25), IN3 => mem_s_1_25_port, 
                           IN4 => n238, Q => n87);
   U62 : AO22X1 port map( IN1 => n239, IN2 => din(24), IN3 => mem_s_1_24_port, 
                           IN4 => n238, Q => n88);
   U63 : AO22X1 port map( IN1 => n240, IN2 => din(23), IN3 => mem_s_1_23_port, 
                           IN4 => n237, Q => n89);
   U64 : AO22X1 port map( IN1 => n240, IN2 => din(22), IN3 => mem_s_1_22_port, 
                           IN4 => n237, Q => n90);
   U65 : AO22X1 port map( IN1 => n240, IN2 => din(21), IN3 => mem_s_1_21_port, 
                           IN4 => n237, Q => n91);
   U66 : AO22X1 port map( IN1 => n239, IN2 => din(20), IN3 => mem_s_1_20_port, 
                           IN4 => n237, Q => n92);
   U67 : AO22X1 port map( IN1 => n240, IN2 => din(19), IN3 => mem_s_1_19_port, 
                           IN4 => n237, Q => n93);
   U68 : AO22X1 port map( IN1 => n239, IN2 => din(18), IN3 => mem_s_1_18_port, 
                           IN4 => n237, Q => n94);
   U69 : AO22X1 port map( IN1 => n240, IN2 => din(17), IN3 => mem_s_1_17_port, 
                           IN4 => n237, Q => n95);
   U70 : AO22X1 port map( IN1 => n239, IN2 => din(16), IN3 => mem_s_1_16_port, 
                           IN4 => n237, Q => n96);
   U71 : AO22X1 port map( IN1 => n240, IN2 => din(15), IN3 => mem_s_1_15_port, 
                           IN4 => n237, Q => n97);
   U72 : AO22X1 port map( IN1 => n239, IN2 => din(14), IN3 => mem_s_1_14_port, 
                           IN4 => n237, Q => n98);
   U73 : AO22X1 port map( IN1 => n239, IN2 => din(13), IN3 => mem_s_1_13_port, 
                           IN4 => n237, Q => n99);
   U74 : AO22X1 port map( IN1 => n239, IN2 => din(12), IN3 => mem_s_1_12_port, 
                           IN4 => n237, Q => n100);
   U75 : AO22X1 port map( IN1 => n239, IN2 => din(11), IN3 => mem_s_1_11_port, 
                           IN4 => n236, Q => n101);
   U76 : AO22X1 port map( IN1 => n239, IN2 => din(10), IN3 => mem_s_1_10_port, 
                           IN4 => n236, Q => n102);
   U77 : AO22X1 port map( IN1 => n239, IN2 => din(9), IN3 => mem_s_1_9_port, 
                           IN4 => n236, Q => n103);
   U78 : AO22X1 port map( IN1 => n240, IN2 => din(8), IN3 => mem_s_1_8_port, 
                           IN4 => n236, Q => n104);
   U79 : AO22X1 port map( IN1 => n240, IN2 => din(7), IN3 => mem_s_1_7_port, 
                           IN4 => n236, Q => n105);
   U80 : AO22X1 port map( IN1 => n239, IN2 => din(6), IN3 => mem_s_1_6_port, 
                           IN4 => n236, Q => n106);
   U81 : AO22X1 port map( IN1 => n239, IN2 => din(5), IN3 => mem_s_1_5_port, 
                           IN4 => n236, Q => n107);
   U82 : AO22X1 port map( IN1 => n240, IN2 => din(4), IN3 => mem_s_1_4_port, 
                           IN4 => n236, Q => n108);
   U83 : AO22X1 port map( IN1 => n240, IN2 => din(3), IN3 => mem_s_1_3_port, 
                           IN4 => n236, Q => n109);
   U84 : AO22X1 port map( IN1 => n240, IN2 => din(2), IN3 => mem_s_1_2_port, 
                           IN4 => n236, Q => n110);
   U85 : AO22X1 port map( IN1 => n240, IN2 => din(1), IN3 => mem_s_1_1_port, 
                           IN4 => n236, Q => n111);
   U86 : AO22X1 port map( IN1 => n240, IN2 => din(0), IN3 => mem_s_1_0_port, 
                           IN4 => n236, Q => n112);
   U87 : AO22X1 port map( IN1 => n235, IN2 => din(31), IN3 => mem_s_2_31_port, 
                           IN4 => n233, Q => n113);
   U88 : AO22X1 port map( IN1 => n235, IN2 => din(30), IN3 => mem_s_2_30_port, 
                           IN4 => n233, Q => n114);
   U89 : AO22X1 port map( IN1 => n235, IN2 => din(29), IN3 => mem_s_2_29_port, 
                           IN4 => n233, Q => n115);
   U90 : AO22X1 port map( IN1 => n235, IN2 => din(28), IN3 => mem_s_2_28_port, 
                           IN4 => n233, Q => n116);
   U91 : AO22X1 port map( IN1 => n234, IN2 => din(27), IN3 => mem_s_2_27_port, 
                           IN4 => n233, Q => n117);
   U92 : AO22X1 port map( IN1 => n234, IN2 => din(26), IN3 => mem_s_2_26_port, 
                           IN4 => n233, Q => n118);
   U93 : AO22X1 port map( IN1 => n234, IN2 => din(25), IN3 => mem_s_2_25_port, 
                           IN4 => n233, Q => n119);
   U94 : AO22X1 port map( IN1 => n234, IN2 => din(24), IN3 => mem_s_2_24_port, 
                           IN4 => n233, Q => n120);
   U95 : AO22X1 port map( IN1 => n235, IN2 => din(23), IN3 => mem_s_2_23_port, 
                           IN4 => n232, Q => n121);
   U96 : AO22X1 port map( IN1 => n235, IN2 => din(22), IN3 => mem_s_2_22_port, 
                           IN4 => n232, Q => n122);
   U97 : AO22X1 port map( IN1 => n235, IN2 => din(21), IN3 => mem_s_2_21_port, 
                           IN4 => n232, Q => n123);
   U98 : AO22X1 port map( IN1 => n234, IN2 => din(20), IN3 => mem_s_2_20_port, 
                           IN4 => n232, Q => n124);
   U99 : AO22X1 port map( IN1 => n235, IN2 => din(19), IN3 => mem_s_2_19_port, 
                           IN4 => n232, Q => n125);
   U100 : AO22X1 port map( IN1 => n234, IN2 => din(18), IN3 => mem_s_2_18_port,
                           IN4 => n232, Q => n126);
   U101 : AO22X1 port map( IN1 => n235, IN2 => din(17), IN3 => mem_s_2_17_port,
                           IN4 => n232, Q => n127);
   U102 : AO22X1 port map( IN1 => n234, IN2 => din(16), IN3 => mem_s_2_16_port,
                           IN4 => n232, Q => n128);
   U103 : AO22X1 port map( IN1 => n235, IN2 => din(15), IN3 => mem_s_2_15_port,
                           IN4 => n232, Q => n129);
   U104 : AO22X1 port map( IN1 => n234, IN2 => din(14), IN3 => mem_s_2_14_port,
                           IN4 => n232, Q => n130);
   U105 : AO22X1 port map( IN1 => n234, IN2 => din(13), IN3 => mem_s_2_13_port,
                           IN4 => n232, Q => n131);
   U106 : AO22X1 port map( IN1 => n234, IN2 => din(12), IN3 => mem_s_2_12_port,
                           IN4 => n232, Q => n132);
   U107 : AO22X1 port map( IN1 => n234, IN2 => din(11), IN3 => mem_s_2_11_port,
                           IN4 => n231, Q => n133);
   U108 : AO22X1 port map( IN1 => n234, IN2 => din(10), IN3 => mem_s_2_10_port,
                           IN4 => n231, Q => n134);
   U109 : AO22X1 port map( IN1 => n234, IN2 => din(9), IN3 => mem_s_2_9_port, 
                           IN4 => n231, Q => n135);
   U110 : AO22X1 port map( IN1 => n235, IN2 => din(8), IN3 => mem_s_2_8_port, 
                           IN4 => n231, Q => n136);
   U111 : AO22X1 port map( IN1 => n235, IN2 => din(7), IN3 => mem_s_2_7_port, 
                           IN4 => n231, Q => n137);
   U112 : AO22X1 port map( IN1 => n234, IN2 => din(6), IN3 => mem_s_2_6_port, 
                           IN4 => n231, Q => n138);
   U113 : AO22X1 port map( IN1 => n234, IN2 => din(5), IN3 => mem_s_2_5_port, 
                           IN4 => n231, Q => n139);
   U114 : AO22X1 port map( IN1 => n235, IN2 => din(4), IN3 => mem_s_2_4_port, 
                           IN4 => n231, Q => n140);
   U115 : AO22X1 port map( IN1 => n235, IN2 => din(3), IN3 => mem_s_2_3_port, 
                           IN4 => n231, Q => n141);
   U116 : AO22X1 port map( IN1 => n235, IN2 => din(2), IN3 => mem_s_2_2_port, 
                           IN4 => n231, Q => n142);
   U117 : AO22X1 port map( IN1 => n235, IN2 => din(1), IN3 => mem_s_2_1_port, 
                           IN4 => n231, Q => n143);
   U118 : AO22X1 port map( IN1 => n235, IN2 => din(0), IN3 => mem_s_2_0_port, 
                           IN4 => n231, Q => n144);
   U119 : NAND3X0 port map( IN1 => n249, IN2 => n25, IN3 => wr_ptr_s_1_port, QN
                           => n28);
   U120 : AO22X1 port map( IN1 => n230, IN2 => din(31), IN3 => mem_s_3_31_port,
                           IN4 => n228, Q => n145);
   U121 : AO22X1 port map( IN1 => n230, IN2 => din(30), IN3 => mem_s_3_30_port,
                           IN4 => n228, Q => n146);
   U122 : AO22X1 port map( IN1 => n230, IN2 => din(29), IN3 => mem_s_3_29_port,
                           IN4 => n228, Q => n147);
   U123 : AO22X1 port map( IN1 => n230, IN2 => din(28), IN3 => mem_s_3_28_port,
                           IN4 => n228, Q => n148);
   U124 : AO22X1 port map( IN1 => n229, IN2 => din(27), IN3 => mem_s_3_27_port,
                           IN4 => n228, Q => n149);
   U125 : AO22X1 port map( IN1 => n229, IN2 => din(26), IN3 => mem_s_3_26_port,
                           IN4 => n228, Q => n150);
   U126 : AO22X1 port map( IN1 => n229, IN2 => din(25), IN3 => mem_s_3_25_port,
                           IN4 => n228, Q => n151);
   U127 : AO22X1 port map( IN1 => n229, IN2 => din(24), IN3 => mem_s_3_24_port,
                           IN4 => n228, Q => n152);
   U128 : AO22X1 port map( IN1 => n230, IN2 => din(23), IN3 => mem_s_3_23_port,
                           IN4 => n227, Q => n153);
   U129 : AO22X1 port map( IN1 => n230, IN2 => din(22), IN3 => mem_s_3_22_port,
                           IN4 => n227, Q => n154);
   U130 : AO22X1 port map( IN1 => n230, IN2 => din(21), IN3 => mem_s_3_21_port,
                           IN4 => n227, Q => n155);
   U131 : AO22X1 port map( IN1 => n229, IN2 => din(20), IN3 => mem_s_3_20_port,
                           IN4 => n227, Q => n156);
   U132 : AO22X1 port map( IN1 => n230, IN2 => din(19), IN3 => mem_s_3_19_port,
                           IN4 => n227, Q => n157);
   U133 : AO22X1 port map( IN1 => n229, IN2 => din(18), IN3 => mem_s_3_18_port,
                           IN4 => n227, Q => n158);
   U134 : AO22X1 port map( IN1 => n230, IN2 => din(17), IN3 => mem_s_3_17_port,
                           IN4 => n227, Q => n159);
   U135 : AO22X1 port map( IN1 => n229, IN2 => din(16), IN3 => mem_s_3_16_port,
                           IN4 => n227, Q => n160);
   U136 : AO22X1 port map( IN1 => n230, IN2 => din(15), IN3 => mem_s_3_15_port,
                           IN4 => n227, Q => n161);
   U137 : AO22X1 port map( IN1 => n229, IN2 => din(14), IN3 => mem_s_3_14_port,
                           IN4 => n227, Q => n162);
   U138 : AO22X1 port map( IN1 => n229, IN2 => din(13), IN3 => mem_s_3_13_port,
                           IN4 => n227, Q => n163);
   U139 : AO22X1 port map( IN1 => n229, IN2 => din(12), IN3 => mem_s_3_12_port,
                           IN4 => n227, Q => n164);
   U140 : AO22X1 port map( IN1 => n229, IN2 => din(11), IN3 => mem_s_3_11_port,
                           IN4 => n226, Q => n165);
   U141 : AO22X1 port map( IN1 => n229, IN2 => din(10), IN3 => mem_s_3_10_port,
                           IN4 => n226, Q => n166);
   U142 : AO22X1 port map( IN1 => n229, IN2 => din(9), IN3 => mem_s_3_9_port, 
                           IN4 => n226, Q => n167);
   U143 : AO22X1 port map( IN1 => n230, IN2 => din(8), IN3 => mem_s_3_8_port, 
                           IN4 => n226, Q => n168);
   U144 : AO22X1 port map( IN1 => n230, IN2 => din(7), IN3 => mem_s_3_7_port, 
                           IN4 => n226, Q => n169);
   U145 : AO22X1 port map( IN1 => n229, IN2 => din(6), IN3 => mem_s_3_6_port, 
                           IN4 => n226, Q => n170);
   U146 : AO22X1 port map( IN1 => n229, IN2 => din(5), IN3 => mem_s_3_5_port, 
                           IN4 => n226, Q => n171);
   U147 : AO22X1 port map( IN1 => n230, IN2 => din(4), IN3 => mem_s_3_4_port, 
                           IN4 => n226, Q => n172);
   U148 : AO22X1 port map( IN1 => n230, IN2 => din(3), IN3 => mem_s_3_3_port, 
                           IN4 => n226, Q => n173);
   U149 : AO22X1 port map( IN1 => n230, IN2 => din(2), IN3 => mem_s_3_2_port, 
                           IN4 => n226, Q => n174);
   U150 : AO22X1 port map( IN1 => n230, IN2 => din(1), IN3 => mem_s_3_1_port, 
                           IN4 => n226, Q => n175);
   U151 : AO22X1 port map( IN1 => n230, IN2 => din(0), IN3 => mem_s_3_0_port, 
                           IN4 => n226, Q => n176);
   U152 : NAND4X0 port map( IN1 => wr_ptr_s_1_port, IN2 => wr_ptr_s_0_port, IN3
                           => n249, IN4 => n251, QN => n29);
   U153 : AO22X1 port map( IN1 => n250, IN2 => wr_ptr_s_0_port, IN3 => n25, IN4
                           => n31, Q => n177);
   U154 : AO22X1 port map( IN1 => n27, IN2 => n31, IN3 => wr_ptr_s_1_port, IN4 
                           => n32, Q => n178);
   U155 : OR2X1 port map( IN1 => n250, IN2 => n25, Q => n32);
   U156 : AND3X1 port map( IN1 => n251, IN2 => n13, IN3 => wr_ptr_s_0_port, Q 
                           => n27);
   U157 : AO22X1 port map( IN1 => N12, IN2 => n33, IN3 => n251, IN4 => n34, Q 
                           => n179);
   U158 : OAI22X1 port map( IN1 => din_ready_port, IN2 => n22, IN3 => n35, IN4 
                           => n21, QN => n34);
   U159 : OA21X1 port map( IN1 => n22, IN2 => n36, IN3 => din_ready_port, Q => 
                           n35);
   U160 : AO22X1 port map( IN1 => entries_s_1_port, IN2 => n33, IN3 => n37, IN4
                           => n251, Q => n180);
   U161 : NAND3X0 port map( IN1 => n40, IN2 => n21, IN3 => n41, QN => n39);
   U162 : XOR2X1 port map( IN1 => n22, IN2 => n248, Q => n41);
   U163 : NAND3X0 port map( IN1 => entries_s_0_port, IN2 => n36, IN3 => 
                           entries_s_1_port, QN => n38);
   U164 : NAND3X0 port map( IN1 => n22, IN2 => n251, IN3 => n248, QN => n42);
   U165 : AO22X1 port map( IN1 => N10, IN2 => n246, IN3 => n43, IN4 => n44, Q 
                           => n181);
   U166 : AO22X1 port map( IN1 => N11, IN2 => n246, IN3 => n45, IN4 => n251, Q 
                           => n182);
   U167 : AO22X1 port map( IN1 => N11, IN2 => n14, IN3 => n46, IN4 => N10, Q =>
                           n45);
   U168 : AO21X1 port map( IN1 => dout_ready, IN2 => dout_valid_port, IN3 => 
                           rst, Q => n44);
   U169 : AO22X1 port map( IN1 => n247, IN2 => entries_s_0_port, IN3 => n47, 
                           IN4 => n40, Q => n183);
   U170 : NAND3X0 port map( IN1 => n36, IN2 => n251, IN3 => n48, QN => n40);
   U171 : NAND3X0 port map( IN1 => n30, IN2 => dout_valid_port, IN3 => 
                           dout_ready, QN => n48);
   U172 : AO21X1 port map( IN1 => dout_ready, IN2 => dout_valid_port, IN3 => 
                           n30, Q => n36);
   U173 : NAND3X0 port map( IN1 => n22, IN2 => n21, IN3 => din_ready_port, QN 
                           => dout_valid_port);
   U3 : INVX0 port map( INP => n239, ZN => n237);
   U4 : INVX0 port map( INP => n240, ZN => n236);
   U5 : INVX0 port map( INP => n239, ZN => n238);
   U6 : INVX0 port map( INP => n245, ZN => n242);
   U7 : INVX0 port map( INP => n244, ZN => n241);
   U8 : INVX0 port map( INP => n234, ZN => n232);
   U9 : INVX0 port map( INP => n235, ZN => n231);
   U10 : INVX0 port map( INP => n229, ZN => n227);
   U11 : INVX0 port map( INP => n230, ZN => n226);
   U12 : INVX0 port map( INP => n245, ZN => n243);
   U13 : INVX0 port map( INP => n234, ZN => n233);
   U14 : INVX0 port map( INP => n229, ZN => n228);
   U15 : INVX0 port map( INP => n26, ZN => n239);
   U16 : INVX0 port map( INP => n26, ZN => n240);
   U17 : INVX0 port map( INP => n36, ZN => n248);
   U18 : NBUFFX2 port map( INP => n200, Z => n210);
   U19 : NBUFFX2 port map( INP => n200, Z => n209);
   U20 : INVX0 port map( INP => n31, ZN => n250);
   U21 : NBUFFX2 port map( INP => n200, Z => n208);
   U174 : INVX0 port map( INP => n30, ZN => n249);
   U175 : NAND2X1 port map( IN1 => n27, IN2 => n249, QN => n26);
   U176 : INVX0 port map( INP => n29, ZN => n229);
   U177 : INVX0 port map( INP => n29, ZN => n230);
   U178 : INVX0 port map( INP => n28, ZN => n234);
   U179 : INVX0 port map( INP => n28, ZN => n235);
   U180 : INVX0 port map( INP => n24, ZN => n244);
   U181 : INVX0 port map( INP => n24, ZN => n245);
   U182 : NAND2X1 port map( IN1 => n251, IN2 => n30, QN => n31);
   U183 : INVX0 port map( INP => n44, ZN => n246);
   U184 : NBUFFX2 port map( INP => n197, Z => n204);
   U185 : NBUFFX2 port map( INP => n197, Z => n203);
   U186 : NBUFFX2 port map( INP => n201, Z => n213);
   U187 : NBUFFX2 port map( INP => n201, Z => n212);
   U188 : NBUFFX2 port map( INP => n198, Z => n206);
   U189 : NBUFFX2 port map( INP => n198, Z => n207);
   U190 : NBUFFX2 port map( INP => n197, Z => n202);
   U191 : NBUFFX2 port map( INP => n201, Z => n211);
   U192 : NBUFFX2 port map( INP => n198, Z => n205);
   U193 : NAND2X1 port map( IN1 => din_valid, IN2 => din_ready_port, QN => n30)
                           ;
   U194 : NOR2X0 port map( IN1 => rst, IN2 => wr_ptr_s_0_port, QN => n25);
   U195 : NAND2X1 port map( IN1 => n40, IN2 => n42, QN => n33);
   U196 : NOR2X0 port map( IN1 => rst, IN2 => N10, QN => n43);
   U197 : NOR2X0 port map( IN1 => N11, IN2 => n246, QN => n46);
   U198 : NOR2X0 port map( IN1 => rst, IN2 => entries_s_0_port, QN => n47);
   U199 : INVX0 port map( INP => n40, ZN => n247);
   U200 : NAND2X1 port map( IN1 => n38, IN2 => n39, QN => n37);
   U201 : INVX0 port map( INP => rst, ZN => n251);
   U202 : NBUFFX2 port map( INP => clk, Z => n224);
   U203 : NBUFFX2 port map( INP => clk, Z => n223);
   U204 : NBUFFX2 port map( INP => clk, Z => n222);
   U205 : NBUFFX2 port map( INP => clk, Z => n221);
   U206 : NBUFFX2 port map( INP => clk, Z => n220);
   U207 : NBUFFX2 port map( INP => clk, Z => n219);
   U208 : NBUFFX2 port map( INP => clk, Z => n218);
   U209 : NBUFFX2 port map( INP => clk, Z => n217);
   U210 : NBUFFX2 port map( INP => clk, Z => n216);
   U211 : NBUFFX2 port map( INP => clk, Z => n215);
   U212 : NBUFFX2 port map( INP => clk, Z => n214);
   U213 : NBUFFX2 port map( INP => clk, Z => n225);
   U214 : NOR2X0 port map( IN1 => n1, IN2 => N10, QN => n201);
   U215 : NOR2X0 port map( IN1 => n1, IN2 => n14, QN => n200);
   U216 : NOR2X0 port map( IN1 => n14, IN2 => N11, QN => n198);
   U217 : NOR2X0 port map( IN1 => N10, IN2 => N11, QN => n197);
   U218 : AO22X1 port map( IN1 => mem_s_1_0_port, IN2 => n205, IN3 => 
                           mem_s_0_0_port, IN4 => n204, Q => n2);
   U219 : AO221X1 port map( IN1 => mem_s_2_0_port, IN2 => n213, IN3 => 
                           mem_s_3_0_port, IN4 => n210, IN5 => n2, Q => dout(0)
                           );
   U220 : AO22X1 port map( IN1 => mem_s_1_1_port, IN2 => n205, IN3 => 
                           mem_s_0_1_port, IN4 => n204, Q => n3);
   U221 : AO221X1 port map( IN1 => mem_s_2_1_port, IN2 => n213, IN3 => 
                           mem_s_3_1_port, IN4 => n210, IN5 => n3, Q => dout(1)
                           );
   U222 : AO22X1 port map( IN1 => mem_s_1_2_port, IN2 => n205, IN3 => 
                           mem_s_0_2_port, IN4 => n204, Q => n4);
   U223 : AO221X1 port map( IN1 => mem_s_2_2_port, IN2 => n213, IN3 => 
                           mem_s_3_2_port, IN4 => n210, IN5 => n4, Q => dout(2)
                           );
   U224 : AO22X1 port map( IN1 => mem_s_1_3_port, IN2 => n205, IN3 => 
                           mem_s_0_3_port, IN4 => n204, Q => n5);
   U225 : AO221X1 port map( IN1 => mem_s_2_3_port, IN2 => n213, IN3 => 
                           mem_s_3_3_port, IN4 => n210, IN5 => n5, Q => dout(3)
                           );
   U226 : AO22X1 port map( IN1 => mem_s_1_4_port, IN2 => n205, IN3 => 
                           mem_s_0_4_port, IN4 => n204, Q => n6);
   U227 : AO221X1 port map( IN1 => mem_s_2_4_port, IN2 => n213, IN3 => 
                           mem_s_3_4_port, IN4 => n210, IN5 => n6, Q => dout(4)
                           );
   U228 : AO22X1 port map( IN1 => mem_s_1_5_port, IN2 => n205, IN3 => 
                           mem_s_0_5_port, IN4 => n204, Q => n7);
   U229 : AO221X1 port map( IN1 => mem_s_2_5_port, IN2 => n213, IN3 => 
                           mem_s_3_5_port, IN4 => n210, IN5 => n7, Q => dout(5)
                           );
   U230 : AO22X1 port map( IN1 => mem_s_1_6_port, IN2 => n205, IN3 => 
                           mem_s_0_6_port, IN4 => n204, Q => n8);
   U231 : AO221X1 port map( IN1 => mem_s_2_6_port, IN2 => n213, IN3 => 
                           mem_s_3_6_port, IN4 => n210, IN5 => n8, Q => dout(6)
                           );
   U232 : AO22X1 port map( IN1 => mem_s_1_7_port, IN2 => n205, IN3 => 
                           mem_s_0_7_port, IN4 => n204, Q => n9);
   U233 : AO221X1 port map( IN1 => mem_s_2_7_port, IN2 => n213, IN3 => 
                           mem_s_3_7_port, IN4 => n210, IN5 => n9, Q => dout(7)
                           );
   U234 : AO22X1 port map( IN1 => mem_s_1_8_port, IN2 => n206, IN3 => 
                           mem_s_0_8_port, IN4 => n204, Q => n10_port);
   U235 : AO221X1 port map( IN1 => mem_s_2_8_port, IN2 => n213, IN3 => 
                           mem_s_3_8_port, IN4 => n210, IN5 => n10_port, Q => 
                           dout(8));
   U236 : AO22X1 port map( IN1 => mem_s_1_9_port, IN2 => n206, IN3 => 
                           mem_s_0_9_port, IN4 => n204, Q => n11_port);
   U237 : AO221X1 port map( IN1 => mem_s_2_9_port, IN2 => n213, IN3 => 
                           mem_s_3_9_port, IN4 => n210, IN5 => n11_port, Q => 
                           dout(9));
   U238 : AO22X1 port map( IN1 => mem_s_1_10_port, IN2 => n206, IN3 => 
                           mem_s_0_10_port, IN4 => n204, Q => n12_port);
   U239 : AO221X1 port map( IN1 => mem_s_2_10_port, IN2 => n213, IN3 => 
                           mem_s_3_10_port, IN4 => n210, IN5 => n12_port, Q => 
                           dout(10));
   U240 : AO22X1 port map( IN1 => mem_s_1_11_port, IN2 => n206, IN3 => 
                           mem_s_0_11_port, IN4 => n204, Q => n15);
   U241 : AO221X1 port map( IN1 => mem_s_2_11_port, IN2 => n213, IN3 => 
                           mem_s_3_11_port, IN4 => n210, IN5 => n15, Q => 
                           dout(11));
   U242 : AO22X1 port map( IN1 => mem_s_1_12_port, IN2 => n206, IN3 => 
                           mem_s_0_12_port, IN4 => n203, Q => n16);
   U243 : AO221X1 port map( IN1 => mem_s_2_12_port, IN2 => n212, IN3 => 
                           mem_s_3_12_port, IN4 => n209, IN5 => n16, Q => 
                           dout(12));
   U244 : AO22X1 port map( IN1 => mem_s_1_13_port, IN2 => n206, IN3 => 
                           mem_s_0_13_port, IN4 => n203, Q => n17);
   U245 : AO221X1 port map( IN1 => mem_s_2_13_port, IN2 => n212, IN3 => 
                           mem_s_3_13_port, IN4 => n209, IN5 => n17, Q => 
                           dout(13));
   U246 : AO22X1 port map( IN1 => mem_s_1_14_port, IN2 => n206, IN3 => 
                           mem_s_0_14_port, IN4 => n203, Q => n18);
   U247 : AO221X1 port map( IN1 => mem_s_2_14_port, IN2 => n212, IN3 => 
                           mem_s_3_14_port, IN4 => n209, IN5 => n18, Q => 
                           dout(14));
   U248 : AO22X1 port map( IN1 => mem_s_1_15_port, IN2 => n206, IN3 => 
                           mem_s_0_15_port, IN4 => n203, Q => n19);
   U249 : AO221X1 port map( IN1 => mem_s_2_15_port, IN2 => n212, IN3 => 
                           mem_s_3_15_port, IN4 => n209, IN5 => n19, Q => 
                           dout(15));
   U250 : AO22X1 port map( IN1 => mem_s_1_16_port, IN2 => n206, IN3 => 
                           mem_s_0_16_port, IN4 => n203, Q => n20);
   U251 : AO221X1 port map( IN1 => mem_s_2_16_port, IN2 => n212, IN3 => 
                           mem_s_3_16_port, IN4 => n209, IN5 => n20, Q => 
                           dout(16));
   U252 : AO22X1 port map( IN1 => mem_s_1_17_port, IN2 => n206, IN3 => 
                           mem_s_0_17_port, IN4 => n203, Q => n23);
   U253 : AO221X1 port map( IN1 => mem_s_2_17_port, IN2 => n212, IN3 => 
                           mem_s_3_17_port, IN4 => n209, IN5 => n23, Q => 
                           dout(17));
   U254 : AO22X1 port map( IN1 => mem_s_1_18_port, IN2 => n206, IN3 => 
                           mem_s_0_18_port, IN4 => n203, Q => n184);
   U255 : AO221X1 port map( IN1 => mem_s_2_18_port, IN2 => n212, IN3 => 
                           mem_s_3_18_port, IN4 => n209, IN5 => n184, Q => 
                           dout(18));
   U256 : AO22X1 port map( IN1 => mem_s_1_19_port, IN2 => n206, IN3 => 
                           mem_s_0_19_port, IN4 => n203, Q => n185);
   U257 : AO221X1 port map( IN1 => mem_s_2_19_port, IN2 => n212, IN3 => 
                           mem_s_3_19_port, IN4 => n209, IN5 => n185, Q => 
                           dout(19));
   U258 : AO22X1 port map( IN1 => mem_s_1_20_port, IN2 => n207, IN3 => 
                           mem_s_0_20_port, IN4 => n203, Q => n186);
   U259 : AO221X1 port map( IN1 => mem_s_2_20_port, IN2 => n212, IN3 => 
                           mem_s_3_20_port, IN4 => n209, IN5 => n186, Q => 
                           dout(20));
   U260 : AO22X1 port map( IN1 => mem_s_1_21_port, IN2 => n207, IN3 => 
                           mem_s_0_21_port, IN4 => n203, Q => n187);
   U261 : AO221X1 port map( IN1 => mem_s_2_21_port, IN2 => n212, IN3 => 
                           mem_s_3_21_port, IN4 => n209, IN5 => n187, Q => 
                           dout(21));
   U262 : AO22X1 port map( IN1 => mem_s_1_22_port, IN2 => n207, IN3 => 
                           mem_s_0_22_port, IN4 => n203, Q => n188);
   U263 : AO221X1 port map( IN1 => mem_s_2_22_port, IN2 => n212, IN3 => 
                           mem_s_3_22_port, IN4 => n209, IN5 => n188, Q => 
                           dout(22));
   U264 : AO22X1 port map( IN1 => mem_s_1_23_port, IN2 => n207, IN3 => 
                           mem_s_0_23_port, IN4 => n203, Q => n189);
   U265 : AO221X1 port map( IN1 => mem_s_2_23_port, IN2 => n212, IN3 => 
                           mem_s_3_23_port, IN4 => n209, IN5 => n189, Q => 
                           dout(23));
   U266 : AO22X1 port map( IN1 => mem_s_1_24_port, IN2 => n207, IN3 => 
                           mem_s_0_24_port, IN4 => n202, Q => n190);
   U267 : AO221X1 port map( IN1 => mem_s_2_24_port, IN2 => n211, IN3 => 
                           mem_s_3_24_port, IN4 => n208, IN5 => n190, Q => 
                           dout(24));
   U268 : AO22X1 port map( IN1 => mem_s_1_25_port, IN2 => n207, IN3 => 
                           mem_s_0_25_port, IN4 => n202, Q => n191);
   U269 : AO221X1 port map( IN1 => mem_s_2_25_port, IN2 => n211, IN3 => 
                           mem_s_3_25_port, IN4 => n208, IN5 => n191, Q => 
                           dout(25));
   U270 : AO22X1 port map( IN1 => mem_s_1_26_port, IN2 => n207, IN3 => 
                           mem_s_0_26_port, IN4 => n202, Q => n192);
   U271 : AO221X1 port map( IN1 => mem_s_2_26_port, IN2 => n211, IN3 => 
                           mem_s_3_26_port, IN4 => n208, IN5 => n192, Q => 
                           dout(26));
   U272 : AO22X1 port map( IN1 => mem_s_1_27_port, IN2 => n207, IN3 => 
                           mem_s_0_27_port, IN4 => n202, Q => n193);
   U273 : AO221X1 port map( IN1 => mem_s_2_27_port, IN2 => n211, IN3 => 
                           mem_s_3_27_port, IN4 => n208, IN5 => n193, Q => 
                           dout(27));
   U274 : AO22X1 port map( IN1 => mem_s_1_28_port, IN2 => n207, IN3 => 
                           mem_s_0_28_port, IN4 => n202, Q => n194);
   U275 : AO221X1 port map( IN1 => mem_s_2_28_port, IN2 => n211, IN3 => 
                           mem_s_3_28_port, IN4 => n208, IN5 => n194, Q => 
                           dout(28));
   U276 : AO22X1 port map( IN1 => mem_s_1_29_port, IN2 => n207, IN3 => 
                           mem_s_0_29_port, IN4 => n202, Q => n195);
   U277 : AO221X1 port map( IN1 => mem_s_2_29_port, IN2 => n211, IN3 => 
                           mem_s_3_29_port, IN4 => n208, IN5 => n195, Q => 
                           dout(29));
   U278 : AO22X1 port map( IN1 => mem_s_1_30_port, IN2 => n207, IN3 => 
                           mem_s_0_30_port, IN4 => n202, Q => n196);
   U279 : AO221X1 port map( IN1 => mem_s_2_30_port, IN2 => n211, IN3 => 
                           mem_s_3_30_port, IN4 => n208, IN5 => n196, Q => 
                           dout(30));
   U280 : AO22X1 port map( IN1 => mem_s_1_31_port, IN2 => n207, IN3 => 
                           mem_s_0_31_port, IN4 => n202, Q => n199);
   U281 : AO221X1 port map( IN1 => mem_s_2_31_port, IN2 => n211, IN3 => 
                           mem_s_3_31_port, IN4 => n208, IN5 => n199, Q => 
                           dout(31));

end SYN_structure;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_LWC_1.all;

entity PostProcessor_1 is

   port( clk, rst : in std_logic;  bdo : in std_logic_vector (31 downto 0);  
         bdo_valid : in std_logic;  bdo_ready : out std_logic;  end_of_block : 
         in std_logic;  bdo_type, bdo_valid_bytes : in std_logic_vector (3 
         downto 0);  msg_auth : in std_logic;  msg_auth_ready : out std_logic; 
         msg_auth_valid : in std_logic;  cmd : in std_logic_vector (31 downto 
         0);  cmd_valid : in std_logic;  cmd_ready : out std_logic;  do_data : 
         out std_logic_vector (31 downto 0);  do_valid, do_last : out std_logic
         ;  do_ready : in std_logic);

end PostProcessor_1;

architecture SYN_PostProcessor of PostProcessor_1 is

   component AND4X1
      port( IN1, IN2, IN3, IN4 : in std_logic;  Q : out std_logic);
   end component;
   
   component NOR4X0
      port( IN1, IN2, IN3, IN4 : in std_logic;  QN : out std_logic);
   end component;
   
   component NOR3X0
      port( IN1, IN2, IN3 : in std_logic;  QN : out std_logic);
   end component;
   
   component OA21X1
      port( IN1, IN2, IN3 : in std_logic;  Q : out std_logic);
   end component;
   
   component AND2X1
      port( IN1, IN2 : in std_logic;  Q : out std_logic);
   end component;
   
   component NAND2X1
      port( IN1, IN2 : in std_logic;  QN : out std_logic);
   end component;
   
   component INVX0
      port( INP : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2X0
      port( IN1, IN2 : in std_logic;  QN : out std_logic);
   end component;
   
   component NAND2X0
      port( IN1, IN2 : in std_logic;  QN : out std_logic);
   end component;
   
   component AND2X4
      port( IN1, IN2 : in std_logic;  Q : out std_logic);
   end component;
   
   component AND2X2
      port( IN1, IN2 : in std_logic;  Q : out std_logic);
   end component;
   
   component DATA_SIPO_1
      port( clk, rst, end_of_input : in std_logic;  data_p : out 
            std_logic_vector (31 downto 0);  data_valid_p : out std_logic;  
            data_ready_p : in std_logic;  data_s : in std_logic_vector (31 
            downto 0);  data_valid_s : in std_logic;  data_ready_s : out 
            std_logic);
   end component;
   
   component StepDownCountLd_N16_step4_1_1
      port( clk, len, ena : in std_logic;  load : in std_logic_vector (15 
            downto 0);  count : out std_logic_vector (15 downto 0));
   end component;
   
   component NAND3X0
      port( IN1, IN2, IN3 : in std_logic;  QN : out std_logic);
   end component;
   
   component AO21X1
      port( IN1, IN2, IN3 : in std_logic;  Q : out std_logic);
   end component;
   
   component NAND4X0
      port( IN1, IN2, IN3, IN4 : in std_logic;  QN : out std_logic);
   end component;
   
   component AO22X1
      port( IN1, IN2, IN3, IN4 : in std_logic;  Q : out std_logic);
   end component;
   
   component AO221X1
      port( IN1, IN2, IN3, IN4, IN5 : in std_logic;  Q : out std_logic);
   end component;
   
   component AND3X1
      port( IN1, IN2, IN3 : in std_logic;  Q : out std_logic);
   end component;
   
   component OA22X1
      port( IN1, IN2, IN3, IN4 : in std_logic;  Q : out std_logic);
   end component;
   
   component OR2X1
      port( IN1, IN2 : in std_logic;  Q : out std_logic);
   end component;
   
   component OR4X1
      port( IN1, IN2, IN3, IN4 : in std_logic;  Q : out std_logic);
   end component;
   
   component AOI222X1
      port( IN1, IN2, IN3, IN4, IN5, IN6 : in std_logic;  QN : out std_logic);
   end component;
   
   component AO222X1
      port( IN1, IN2, IN3, IN4, IN5, IN6 : in std_logic;  Q : out std_logic);
   end component;
   
   component OA221X1
      port( IN1, IN2, IN3, IN4, IN5 : in std_logic;  Q : out std_logic);
   end component;
   
   component DFFX1
      port( D, CLK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFSSRX1
      port( D, RSTB, SETB, CLK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal do_valid_port, do_last_port, bdo_cleared_31_port, bdo_cleared_30_port
      , bdo_cleared_29_port, bdo_cleared_28_port, bdo_cleared_27_port, 
      bdo_cleared_26_port, bdo_cleared_25_port, bdo_cleared_24_port, 
      bdo_cleared_23_port, bdo_cleared_22_port, bdo_cleared_21_port, 
      bdo_cleared_20_port, bdo_cleared_19_port, bdo_cleared_18_port, 
      bdo_cleared_17_port, bdo_cleared_16_port, bdo_cleared_15_port, 
      bdo_cleared_14_port, bdo_cleared_13_port, bdo_cleared_12_port, 
      bdo_cleared_11_port, bdo_cleared_10_port, bdo_cleared_9_port, 
      bdo_cleared_8_port, bdo_cleared_7_port, bdo_cleared_6_port, 
      bdo_cleared_5_port, bdo_cleared_4_port, bdo_cleared_3_port, 
      bdo_cleared_2_port, bdo_cleared_1_port, bdo_cleared_0_port, en_SegLenCnt,
      dout_SegLenCnt_15_port, dout_SegLenCnt_14_port, dout_SegLenCnt_13_port, 
      dout_SegLenCnt_12_port, dout_SegLenCnt_11_port, dout_SegLenCnt_10_port, 
      dout_SegLenCnt_9_port, dout_SegLenCnt_8_port, dout_SegLenCnt_7_port, 
      dout_SegLenCnt_6_port, dout_SegLenCnt_5_port, dout_SegLenCnt_4_port, 
      dout_SegLenCnt_3_port, dout_SegLenCnt_2_port, dout_SegLenCnt_1_port, 
      dout_SegLenCnt_0_port, N40, eot, decrypt, bdo_ready_p, bdo_valid_p, 
      bdo_p_31_port, bdo_p_30_port, bdo_p_29_port, bdo_p_28_port, bdo_p_27_port
      , bdo_p_26_port, bdo_p_25_port, bdo_p_24_port, bdo_p_23_port, 
      bdo_p_22_port, bdo_p_21_port, bdo_p_20_port, bdo_p_19_port, bdo_p_18_port
      , bdo_p_17_port, bdo_p_16_port, bdo_p_15_port, bdo_p_14_port, 
      bdo_p_13_port, bdo_p_12_port, bdo_p_11_port, bdo_p_10_port, bdo_p_9_port,
      bdo_p_8_port, bdo_p_7_port, bdo_p_6_port, bdo_p_5_port, bdo_p_4_port, 
      bdo_p_3_port, bdo_p_2_port, bdo_p_1_port, bdo_p_0_port, pr_state_3_port, 
      pr_state_2_port, pr_state_1_port, pr_state_0_port, n7, n8, n21, n22, n26,
      n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40_port
      , n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, 
      n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69
      , n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, 
      n84, n85, n86, n87, n1, n2, n3, n4, n5, n6, n9, n10, n11, n12, n13, n14, 
      n15, n16, n17, n18, n19, msg_auth_ready_port, n23, n24, n25, n88, n_3220,
      n_3221 : std_logic;

begin
   msg_auth_ready <= msg_auth_ready_port;
   do_valid <= do_valid_port;
   do_last <= do_last_port;
   
   pr_state_reg_0_inst : DFFX1 port map( D => n87, CLK => clk, Q => 
                           pr_state_0_port, QN => n22);
   pr_state_reg_2_inst : DFFX1 port map( D => n86, CLK => clk, Q => 
                           pr_state_2_port, QN => n21);
   eot_reg : DFFX1 port map( D => n83, CLK => clk, Q => eot, QN => n7);
   pr_state_reg_1_inst : DFFX1 port map( D => n85, CLK => clk, Q => 
                           pr_state_1_port, QN => n_3220);
   pr_state_reg_3_inst : DFFSSRX1 port map( D => n54, RSTB => n25, SETB => n24,
                           CLK => clk, Q => pr_state_3_port, QN => n_3221);
   decrypt_reg : DFFX1 port map( D => n84, CLK => clk, Q => decrypt, QN => n8);
   U45 : AO22X1 port map( IN1 => cmd(25), IN2 => n14, IN3 => eot, IN4 => n26, Q
                           => n83);
   U46 : NAND4X0 port map( IN1 => n15, IN2 => n27, IN3 => n28, IN4 => n29, QN 
                           => n26);
   U47 : NOR3X0 port map( IN1 => n30, IN2 => do_last_port, IN3 => n31, QN => 
                           n29);
   U48 : AO22X1 port map( IN1 => cmd(28), IN2 => n10, IN3 => decrypt, IN4 => 
                           n32, Q => n84);
   U49 : NAND4X0 port map( IN1 => n28, IN2 => n15, IN3 => cmd_valid, IN4 => n33
                           , QN => n32);
   U50 : AO22X1 port map( IN1 => n34, IN2 => pr_state_1_port, IN3 => n35, IN4 
                           => n25, Q => n85);
   U51 : NAND4X0 port map( IN1 => n36, IN2 => n37, IN3 => n38, IN4 => n39, QN 
                           => n35);
   U52 : OA221X1 port map( IN1 => n40_port, IN2 => n18, IN3 => n15, IN4 => n88,
                           IN5 => n41, Q => n39);
   U53 : NAND3X0 port map( IN1 => cmd_valid, IN2 => n44, IN3 => n30, QN => n37)
                           ;
   U54 : NAND3X0 port map( IN1 => cmd(31), IN2 => n12, IN3 => n45, QN => n44);
   U55 : NAND3X0 port map( IN1 => en_SegLenCnt, IN2 => n7, IN3 => N40, QN => 
                           n36);
   U56 : AO22X1 port map( IN1 => n34, IN2 => pr_state_2_port, IN3 => n46, IN4 
                           => n25, Q => n86);
   U57 : NAND4X0 port map( IN1 => n47, IN2 => n48, IN3 => n49, IN4 => n50, QN 
                           => n46);
   U58 : OA22X1 port map( IN1 => n40_port, IN2 => n51, IN3 => msg_auth_valid, 
                           IN4 => n27, Q => n50);
   U59 : NAND4X0 port map( IN1 => N40, IN2 => bdo_valid_p, IN3 => do_ready, IN4
                           => n7, QN => n53);
   U60 : AO222X1 port map( IN1 => msg_auth_valid, IN2 => msg_auth_ready_port, 
                           IN3 => n40_port, IN4 => n42, IN5 => pr_state_3_port,
                           IN6 => n88, Q => n54);
   U61 : AO22X1 port map( IN1 => n34, IN2 => pr_state_0_port, IN3 => n55, IN4 
                           => n25, Q => n87);
   U62 : NAND4X0 port map( IN1 => n41, IN2 => n56, IN3 => n9, IN4 => n57, QN =>
                           n55);
   U63 : AOI222X1 port map( IN1 => cmd_valid, IN2 => n30, IN3 => n88, IN4 => 
                           n58, IN5 => n42, IN6 => n40_port, QN => n57);
   U64 : AND3X1 port map( IN1 => bdo_valid_p, IN2 => do_ready, IN3 => 
                           end_of_block, Q => n40_port);
   U65 : AO21X1 port map( IN1 => N40, IN2 => en_SegLenCnt, IN3 => n59, Q => n43
                           );
   U66 : OR4X1 port map( IN1 => n64, IN2 => cmd(0), IN3 => cmd(10), IN4 => 
                           cmd(11), Q => n63);
   U67 : OR4X1 port map( IN1 => cmd(12), IN2 => cmd(13), IN3 => cmd(14), IN4 =>
                           cmd(15), Q => n62);
   U68 : OR4X1 port map( IN1 => cmd(1), IN2 => cmd(2), IN3 => cmd(3), IN4 => 
                           cmd(4), Q => n61);
   U69 : OR4X1 port map( IN1 => cmd(5), IN2 => cmd(6), IN3 => n65, IN4 => 
                           cmd(7), Q => n60);
   U70 : OR2X1 port map( IN1 => cmd(9), IN2 => cmd(8), Q => n65);
   U71 : OA22X1 port map( IN1 => n27, IN2 => msg_auth_valid, IN3 => n64, IN4 =>
                           n66, Q => n41);
   U72 : AND2X1 port map( IN1 => do_ready, IN2 => cmd_valid, Q => n66);
   U73 : AND2X1 port map( IN1 => n31, IN2 => n25, Q => n34);
   U74 : OA21X1 port map( IN1 => pr_state_2_port, IN2 => pr_state_1_port, IN3 
                           => pr_state_3_port, Q => n31);
   U75 : NAND3X0 port map( IN1 => n67, IN2 => pr_state_0_port, IN3 => 
                           pr_state_1_port, QN => n27);
   U76 : NAND3X0 port map( IN1 => do_ready, IN2 => cmd_valid, IN3 => n23, QN =>
                           n48);
   U77 : AND3X1 port map( IN1 => n52, IN2 => do_ready, IN3 => bdo_valid_p, Q =>
                           en_SegLenCnt);
   U78 : AO22X1 port map( IN1 => bdo_p_9_port, IN2 => n68, IN3 => cmd(9), IN4 
                           => n6, Q => do_data(9));
   U79 : AO22X1 port map( IN1 => bdo_p_8_port, IN2 => n68, IN3 => cmd(8), IN4 
                           => n6, Q => do_data(8));
   U80 : AO22X1 port map( IN1 => bdo_p_7_port, IN2 => n68, IN3 => cmd(7), IN4 
                           => n6, Q => do_data(7));
   U81 : AO22X1 port map( IN1 => bdo_p_6_port, IN2 => n68, IN3 => cmd(6), IN4 
                           => n6, Q => do_data(6));
   U82 : AO221X1 port map( IN1 => cmd(5), IN2 => n6, IN3 => bdo_p_5_port, IN4 
                           => n68, IN5 => n13, Q => do_data(5));
   U83 : AO221X1 port map( IN1 => cmd(4), IN2 => n6, IN3 => bdo_p_4_port, IN4 
                           => n68, IN5 => n16, Q => do_data(4));
   U84 : AO22X1 port map( IN1 => bdo_p_3_port, IN2 => n68, IN3 => cmd(3), IN4 
                           => n6, Q => do_data(3));
   U85 : NAND3X0 port map( IN1 => n70, IN2 => n17, IN3 => n15, QN => 
                           do_data(31));
   U86 : NAND3X0 port map( IN1 => n71, IN2 => n17, IN3 => n72, QN => 
                           do_data(30));
   U87 : AO22X1 port map( IN1 => bdo_p_2_port, IN2 => n68, IN3 => cmd(2), IN4 
                           => n6, Q => do_data(2));
   U88 : AO21X1 port map( IN1 => bdo_p_29_port, IN2 => n68, IN3 => do_last_port
                           , Q => do_data(29));
   U89 : AO221X1 port map( IN1 => n6, IN2 => n8, IN3 => bdo_p_28_port, IN4 => 
                           n68, IN5 => n73, Q => do_data(28));
   U90 : AND2X1 port map( IN1 => bdo_p_27_port, IN2 => n68, Q => do_data(27));
   U91 : AND2X1 port map( IN1 => bdo_p_26_port, IN2 => n68, Q => do_data(26));
   U92 : AO221X1 port map( IN1 => n6, IN2 => cmd(25), IN3 => bdo_p_25_port, IN4
                           => n68, IN5 => n75, Q => do_data(25));
   U93 : AO221X1 port map( IN1 => n76, IN2 => n6, IN3 => bdo_p_24_port, IN4 => 
                           n68, IN5 => n75, Q => do_data(24));
   U94 : AND2X1 port map( IN1 => cmd(25), IN2 => decrypt, Q => n76);
   U95 : AND2X1 port map( IN1 => bdo_p_23_port, IN2 => n68, Q => do_data(23));
   U96 : AND2X1 port map( IN1 => bdo_p_22_port, IN2 => n68, Q => do_data(22));
   U97 : AND2X1 port map( IN1 => bdo_p_21_port, IN2 => n68, Q => do_data(21));
   U98 : AND2X1 port map( IN1 => bdo_p_20_port, IN2 => n68, Q => do_data(20));
   U99 : AO22X1 port map( IN1 => bdo_p_1_port, IN2 => n68, IN3 => cmd(1), IN4 
                           => n6, Q => do_data(1));
   U100 : AND2X1 port map( IN1 => bdo_p_19_port, IN2 => n68, Q => do_data(19));
   U101 : AND2X1 port map( IN1 => bdo_p_18_port, IN2 => n68, Q => do_data(18));
   U102 : AND2X1 port map( IN1 => bdo_p_17_port, IN2 => n68, Q => do_data(17));
   U103 : AND2X1 port map( IN1 => bdo_p_16_port, IN2 => n68, Q => do_data(16));
   U104 : AO22X1 port map( IN1 => bdo_p_15_port, IN2 => n68, IN3 => cmd(15), 
                           IN4 => n6, Q => do_data(15));
   U105 : AO22X1 port map( IN1 => bdo_p_14_port, IN2 => n68, IN3 => cmd(14), 
                           IN4 => n6, Q => do_data(14));
   U106 : AO22X1 port map( IN1 => bdo_p_13_port, IN2 => n68, IN3 => cmd(13), 
                           IN4 => n6, Q => do_data(13));
   U107 : AO22X1 port map( IN1 => bdo_p_12_port, IN2 => n68, IN3 => cmd(12), 
                           IN4 => n6, Q => do_data(12));
   U108 : AO22X1 port map( IN1 => bdo_p_11_port, IN2 => n68, IN3 => cmd(11), 
                           IN4 => n6, Q => do_data(11));
   U109 : AO22X1 port map( IN1 => bdo_p_10_port, IN2 => n68, IN3 => cmd(10), 
                           IN4 => n6, Q => do_data(10));
   U110 : AO22X1 port map( IN1 => bdo_p_0_port, IN2 => n68, IN3 => cmd(0), IN4 
                           => n6, Q => do_data(0));
   U111 : AND2X1 port map( IN1 => do_valid_port, IN2 => n19, Q => n68);
   U112 : NAND4X0 port map( IN1 => n15, IN2 => n77, IN3 => n78, IN4 => n17, QN 
                           => do_valid_port);
   U113 : NAND3X0 port map( IN1 => pr_state_3_port, IN2 => n21, IN3 => n58, QN 
                           => n79);
   U114 : NAND3X0 port map( IN1 => pr_state_3_port, IN2 => n21, IN3 => n80, QN 
                           => n74);
   U115 : AO21X1 port map( IN1 => n23, IN2 => do_ready, IN3 => n30, Q => 
                           cmd_ready);
   U116 : AND2X1 port map( IN1 => n81, IN2 => n80, Q => n30);
   U117 : NAND3X0 port map( IN1 => pr_state_0_port, IN2 => n81, IN3 => 
                           pr_state_1_port, QN => n64);
   U118 : AND2X1 port map( IN1 => n67, IN2 => n80, Q => n52);
   U119 : NAND3X0 port map( IN1 => n81, IN2 => n22, IN3 => pr_state_1_port, QN 
                           => n82);
   U120 : NAND3X0 port map( IN1 => n67, IN2 => n22, IN3 => pr_state_1_port, QN 
                           => n51);
   U121 : AND2X1 port map( IN1 => bdo_valid_bytes(1), IN2 => bdo(9), Q => 
                           bdo_cleared_9_port);
   U122 : AND2X1 port map( IN1 => bdo(8), IN2 => bdo_valid_bytes(1), Q => 
                           bdo_cleared_8_port);
   U123 : AND2X1 port map( IN1 => bdo_valid_bytes(0), IN2 => bdo(7), Q => 
                           bdo_cleared_7_port);
   U125 : AND2X1 port map( IN1 => bdo(5), IN2 => bdo_valid_bytes(0), Q => 
                           bdo_cleared_5_port);
   U126 : AND2X1 port map( IN1 => bdo(4), IN2 => bdo_valid_bytes(0), Q => 
                           bdo_cleared_4_port);
   U127 : AND2X1 port map( IN1 => bdo(3), IN2 => bdo_valid_bytes(0), Q => 
                           bdo_cleared_3_port);
   U128 : AND2X1 port map( IN1 => bdo_valid_bytes(3), IN2 => bdo(31), Q => 
                           bdo_cleared_31_port);
   U135 : AND2X1 port map( IN1 => bdo(25), IN2 => bdo_valid_bytes(3), Q => 
                           bdo_cleared_25_port);
   U136 : AND2X1 port map( IN1 => bdo(24), IN2 => bdo_valid_bytes(3), Q => 
                           bdo_cleared_24_port);
   U139 : AND2X1 port map( IN1 => bdo(21), IN2 => bdo_valid_bytes(2), Q => 
                           bdo_cleared_21_port);
   U140 : AND2X1 port map( IN1 => bdo(20), IN2 => bdo_valid_bytes(2), Q => 
                           bdo_cleared_20_port);
   U141 : AND2X1 port map( IN1 => bdo(1), IN2 => bdo_valid_bytes(0), Q => 
                           bdo_cleared_1_port);
   U142 : AND2X1 port map( IN1 => bdo(19), IN2 => bdo_valid_bytes(2), Q => 
                           bdo_cleared_19_port);
   U143 : AND2X1 port map( IN1 => bdo(18), IN2 => bdo_valid_bytes(2), Q => 
                           bdo_cleared_18_port);
   U145 : AND2X1 port map( IN1 => bdo(16), IN2 => bdo_valid_bytes(2), Q => 
                           bdo_cleared_16_port);
   U146 : AND2X1 port map( IN1 => bdo(15), IN2 => bdo_valid_bytes(1), Q => 
                           bdo_cleared_15_port);
   U147 : AND2X1 port map( IN1 => bdo(14), IN2 => bdo_valid_bytes(1), Q => 
                           bdo_cleared_14_port);
   U148 : AND2X1 port map( IN1 => bdo(13), IN2 => bdo_valid_bytes(1), Q => 
                           bdo_cleared_13_port);
   U151 : AND2X1 port map( IN1 => bdo(10), IN2 => bdo_valid_bytes(1), Q => 
                           bdo_cleared_10_port);
   U152 : AND2X1 port map( IN1 => bdo(0), IN2 => bdo_valid_bytes(0), Q => 
                           bdo_cleared_0_port);
   SegLen : StepDownCountLd_N16_step4_1_1 port map( clk => clk, len => n11, ena
                           => en_SegLenCnt, load(15) => cmd(15), load(14) => 
                           cmd(14), load(13) => cmd(13), load(12) => cmd(12), 
                           load(11) => cmd(11), load(10) => cmd(10), load(9) =>
                           cmd(9), load(8) => cmd(8), load(7) => cmd(7), 
                           load(6) => cmd(6), load(5) => cmd(5), load(4) => 
                           cmd(4), load(3) => cmd(3), load(2) => cmd(2), 
                           load(1) => cmd(1), load(0) => cmd(0), count(15) => 
                           dout_SegLenCnt_15_port, count(14) => 
                           dout_SegLenCnt_14_port, count(13) => 
                           dout_SegLenCnt_13_port, count(12) => 
                           dout_SegLenCnt_12_port, count(11) => 
                           dout_SegLenCnt_11_port, count(10) => 
                           dout_SegLenCnt_10_port, count(9) => 
                           dout_SegLenCnt_9_port, count(8) => 
                           dout_SegLenCnt_8_port, count(7) => 
                           dout_SegLenCnt_7_port, count(6) => 
                           dout_SegLenCnt_6_port, count(5) => 
                           dout_SegLenCnt_5_port, count(4) => 
                           dout_SegLenCnt_4_port, count(3) => 
                           dout_SegLenCnt_3_port, count(2) => 
                           dout_SegLenCnt_2_port, count(1) => 
                           dout_SegLenCnt_1_port, count(0) => 
                           dout_SegLenCnt_0_port);
   bdoSIPO : DATA_SIPO_1 port map( clk => clk, rst => rst, end_of_input => 
                           end_of_block, data_p(31) => bdo_p_31_port, 
                           data_p(30) => bdo_p_30_port, data_p(29) => 
                           bdo_p_29_port, data_p(28) => bdo_p_28_port, 
                           data_p(27) => bdo_p_27_port, data_p(26) => 
                           bdo_p_26_port, data_p(25) => bdo_p_25_port, 
                           data_p(24) => bdo_p_24_port, data_p(23) => 
                           bdo_p_23_port, data_p(22) => bdo_p_22_port, 
                           data_p(21) => bdo_p_21_port, data_p(20) => 
                           bdo_p_20_port, data_p(19) => bdo_p_19_port, 
                           data_p(18) => bdo_p_18_port, data_p(17) => 
                           bdo_p_17_port, data_p(16) => bdo_p_16_port, 
                           data_p(15) => bdo_p_15_port, data_p(14) => 
                           bdo_p_14_port, data_p(13) => bdo_p_13_port, 
                           data_p(12) => bdo_p_12_port, data_p(11) => 
                           bdo_p_11_port, data_p(10) => bdo_p_10_port, 
                           data_p(9) => bdo_p_9_port, data_p(8) => bdo_p_8_port
                           , data_p(7) => bdo_p_7_port, data_p(6) => 
                           bdo_p_6_port, data_p(5) => bdo_p_5_port, data_p(4) 
                           => bdo_p_4_port, data_p(3) => bdo_p_3_port, 
                           data_p(2) => bdo_p_2_port, data_p(1) => bdo_p_1_port
                           , data_p(0) => bdo_p_0_port, data_valid_p => 
                           bdo_valid_p, data_ready_p => bdo_ready_p, data_s(31)
                           => bdo_cleared_31_port, data_s(30) => 
                           bdo_cleared_30_port, data_s(29) => 
                           bdo_cleared_29_port, data_s(28) => 
                           bdo_cleared_28_port, data_s(27) => 
                           bdo_cleared_27_port, data_s(26) => 
                           bdo_cleared_26_port, data_s(25) => 
                           bdo_cleared_25_port, data_s(24) => 
                           bdo_cleared_24_port, data_s(23) => 
                           bdo_cleared_23_port, data_s(22) => 
                           bdo_cleared_22_port, data_s(21) => 
                           bdo_cleared_21_port, data_s(20) => 
                           bdo_cleared_20_port, data_s(19) => 
                           bdo_cleared_19_port, data_s(18) => 
                           bdo_cleared_18_port, data_s(17) => 
                           bdo_cleared_17_port, data_s(16) => 
                           bdo_cleared_16_port, data_s(15) => 
                           bdo_cleared_15_port, data_s(14) => 
                           bdo_cleared_14_port, data_s(13) => 
                           bdo_cleared_13_port, data_s(12) => 
                           bdo_cleared_12_port, data_s(11) => 
                           bdo_cleared_11_port, data_s(10) => 
                           bdo_cleared_10_port, data_s(9) => bdo_cleared_9_port
                           , data_s(8) => bdo_cleared_8_port, data_s(7) => 
                           bdo_cleared_7_port, data_s(6) => bdo_cleared_6_port,
                           data_s(5) => bdo_cleared_5_port, data_s(4) => 
                           bdo_cleared_4_port, data_s(3) => bdo_cleared_3_port,
                           data_s(2) => bdo_cleared_2_port, data_s(1) => 
                           bdo_cleared_1_port, data_s(0) => bdo_cleared_0_port,
                           data_valid_s => bdo_valid, data_ready_s => bdo_ready
                           );
   U3 : AND2X1 port map( IN1 => bdo(2), IN2 => bdo_valid_bytes(0), Q => 
                           bdo_cleared_2_port);
   U4 : AND2X1 port map( IN1 => bdo(6), IN2 => bdo_valid_bytes(0), Q => 
                           bdo_cleared_6_port);
   U5 : AND2X2 port map( IN1 => bdo(22), IN2 => bdo_valid_bytes(2), Q => 
                           bdo_cleared_22_port);
   U6 : AND2X4 port map( IN1 => bdo_valid_bytes(2), IN2 => bdo(23), Q => 
                           bdo_cleared_23_port);
   U7 : AND2X4 port map( IN1 => bdo(27), IN2 => bdo_valid_bytes(3), Q => 
                           bdo_cleared_27_port);
   U8 : AND2X4 port map( IN1 => bdo(26), IN2 => bdo_valid_bytes(3), Q => 
                           bdo_cleared_26_port);
   U9 : AND2X4 port map( IN1 => bdo(12), IN2 => bdo_valid_bytes(1), Q => 
                           bdo_cleared_12_port);
   U10 : NAND2X0 port map( IN1 => n58, IN2 => n81, QN => n69);
   U11 : NAND2X0 port map( IN1 => n67, IN2 => n58, QN => n47);
   U12 : INVX0 port map( INP => n75, ZN => n15);
   U13 : INVX0 port map( INP => n71, ZN => n6);
   U14 : NAND2X1 port map( IN1 => n69, IN2 => n47, QN => n75);
   U15 : INVX0 port map( INP => n34, ZN => n24);
   U16 : NAND2X1 port map( IN1 => n23, IN2 => do_valid_port, QN => n71);
   U17 : INVX0 port map( INP => n28, ZN => n19);
   U18 : NAND2X1 port map( IN1 => bdo_p_31_port, IN2 => n68, QN => n70);
   U19 : NAND2X1 port map( IN1 => bdo_p_30_port, IN2 => n68, QN => n72);
   U20 : AND2X1 port map( IN1 => bdo(30), IN2 => bdo_valid_bytes(3), Q => 
                           bdo_cleared_30_port);
   U21 : AND2X1 port map( IN1 => bdo(17), IN2 => bdo_valid_bytes(2), Q => 
                           bdo_cleared_17_port);
   U22 : NOR2X0 port map( IN1 => n42, IN2 => n52, QN => n28);
   U23 : NOR2X0 port map( IN1 => n28, IN2 => n88, QN => bdo_ready_p);
   U24 : NOR4X0 port map( IN1 => n60, IN2 => n61, IN3 => n62, IN4 => n63, QN =>
                           n59);
   U25 : INVX0 port map( INP => n42, ZN => n18);
   U26 : INVX0 port map( INP => n27, ZN => msg_auth_ready_port);
   U27 : INVX0 port map( INP => n48, ZN => n11);
   U28 : INVX0 port map( INP => n64, ZN => n23);
   U29 : NAND2X1 port map( IN1 => bdo_valid_p, IN2 => n19, QN => n78);
   U30 : NAND2X1 port map( IN1 => n23, IN2 => cmd_valid, QN => n77);
   U31 : INVX0 port map( INP => do_last_port, ZN => n17);
   U32 : INVX0 port map( INP => n47, ZN => n16);
   U33 : INVX0 port map( INP => n69, ZN => n13);
   U34 : AND2X1 port map( IN1 => bdo(11), IN2 => bdo_valid_bytes(1), Q => 
                           bdo_cleared_11_port);
   U35 : AND2X1 port map( IN1 => bdo(29), IN2 => bdo_valid_bytes(3), Q => 
                           bdo_cleared_29_port);
   U36 : NOR2X0 port map( IN1 => n21, IN2 => pr_state_3_port, QN => n67);
   U37 : NOR2X0 port map( IN1 => pr_state_2_port, IN2 => pr_state_3_port, QN =>
                           n81);
   U38 : NAND2X1 port map( IN1 => n51, IN2 => n82, QN => n42);
   U39 : NOR2X0 port map( IN1 => pr_state_0_port, IN2 => pr_state_1_port, QN =>
                           n80);
   U40 : NAND2X1 port map( IN1 => decrypt, IN2 => n43, QN => n38);
   U41 : NAND2X1 port map( IN1 => msg_auth, IN2 => msg_auth_ready_port, QN => 
                           n56);
   U42 : INVX0 port map( INP => n43, ZN => n9);
   U43 : NAND2X0 port map( IN1 => n52, IN2 => n53, QN => n49);
   U44 : NOR2X0 port map( IN1 => n22, IN2 => pr_state_1_port, QN => n58);
   U124 : NAND2X1 port map( IN1 => n74, IN2 => n79, QN => do_last_port);
   U129 : INVX0 port map( INP => cmd(28), ZN => n12);
   U130 : NOR2X0 port map( IN1 => cmd(30), IN2 => cmd(29), QN => n45);
   U131 : INVX0 port map( INP => n26, ZN => n14);
   U132 : INVX0 port map( INP => n32, ZN => n10);
   U133 : NOR4X0 port map( IN1 => do_last_port, IN2 => n31, IN3 => 
                           msg_auth_ready_port, IN4 => n23, QN => n33);
   U134 : INVX0 port map( INP => rst, ZN => n25);
   U137 : INVX0 port map( INP => do_ready, ZN => n88);
   U138 : NAND2X1 port map( IN1 => n69, IN2 => n74, QN => n73);
   U144 : AND2X1 port map( IN1 => bdo(28), IN2 => bdo_valid_bytes(3), Q => 
                           bdo_cleared_28_port);
   U149 : OA21X1 port map( IN1 => dout_SegLenCnt_0_port, IN2 => 
                           dout_SegLenCnt_1_port, IN3 => dout_SegLenCnt_2_port,
                           Q => n1);
   U150 : NOR3X0 port map( IN1 => n1, IN2 => dout_SegLenCnt_11_port, IN3 => 
                           dout_SegLenCnt_10_port, QN => n5);
   U153 : NOR4X0 port map( IN1 => dout_SegLenCnt_15_port, IN2 => 
                           dout_SegLenCnt_14_port, IN3 => 
                           dout_SegLenCnt_13_port, IN4 => 
                           dout_SegLenCnt_12_port, QN => n4);
   U154 : NOR3X0 port map( IN1 => dout_SegLenCnt_3_port, IN2 => 
                           dout_SegLenCnt_5_port, IN3 => dout_SegLenCnt_4_port,
                           QN => n3);
   U155 : NOR4X0 port map( IN1 => dout_SegLenCnt_9_port, IN2 => 
                           dout_SegLenCnt_8_port, IN3 => dout_SegLenCnt_7_port,
                           IN4 => dout_SegLenCnt_6_port, QN => n2);
   U156 : AND4X1 port map( IN1 => n5, IN2 => n4, IN3 => n3, IN4 => n2, Q => N40
                           );

end SYN_PostProcessor;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_LWC_1.all;

entity CryptoCore_1 is

   port( clk, rst : in std_logic;  key : in std_logic_vector (31 downto 0);  
         key_valid : in std_logic;  key_ready : out std_logic;  bdi : in 
         std_logic_vector (31 downto 0);  bdi_valid : in std_logic;  bdi_ready 
         : out std_logic;  bdi_pad_loc, bdi_valid_bytes : in std_logic_vector 
         (3 downto 0);  bdi_size : in std_logic_vector (2 downto 0);  bdi_eot, 
         bdi_eoi : in std_logic;  bdi_type : in std_logic_vector (3 downto 0); 
         decrypt_in, key_update, hash_in : in std_logic;  bdo : out 
         std_logic_vector (31 downto 0);  bdo_valid : out std_logic;  bdo_ready
         : in std_logic;  bdo_type, bdo_valid_bytes : out std_logic_vector (3 
         downto 0);  end_of_block, msg_auth_valid : out std_logic;  
         msg_auth_ready : in std_logic;  msg_auth : out std_logic);

end CryptoCore_1;

architecture SYN_behavioral of CryptoCore_1 is

   component NOR2X0
      port( IN1, IN2 : in std_logic;  QN : out std_logic);
   end component;
   
   component NAND2X0
      port( IN1, IN2 : in std_logic;  QN : out std_logic);
   end component;
   
   component AO21X1
      port( IN1, IN2, IN3 : in std_logic;  Q : out std_logic);
   end component;
   
   component AOI21X1
      port( IN1, IN2, IN3 : in std_logic;  QN : out std_logic);
   end component;
   
   component INVX0
      port( INP : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2X1
      port( IN1, IN2 : in std_logic;  QN : out std_logic);
   end component;
   
   component NAND3X1
      port( IN1, IN2, IN3 : in std_logic;  QN : out std_logic);
   end component;
   
   component NOR3X0
      port( IN1, IN2, IN3 : in std_logic;  QN : out std_logic);
   end component;
   
   component NBUFFX2
      port( INP : in std_logic;  Z : out std_logic);
   end component;
   
   component AO22X1
      port( IN1, IN2, IN3, IN4 : in std_logic;  Q : out std_logic);
   end component;
   
   component NAND3X0
      port( IN1, IN2, IN3 : in std_logic;  QN : out std_logic);
   end component;
   
   component AND4X1
      port( IN1, IN2, IN3, IN4 : in std_logic;  Q : out std_logic);
   end component;
   
   component NOR4X0
      port( IN1, IN2, IN3, IN4 : in std_logic;  QN : out std_logic);
   end component;
   
   component AND2X1
      port( IN1, IN2 : in std_logic;  Q : out std_logic);
   end component;
   
   component NAND4X0
      port( IN1, IN2, IN3, IN4 : in std_logic;  QN : out std_logic);
   end component;
   
   component OR2X1
      port( IN1, IN2 : in std_logic;  Q : out std_logic);
   end component;
   
   component AND3X1
      port( IN1, IN2, IN3 : in std_logic;  Q : out std_logic);
   end component;
   
   component AND2X2
      port( IN1, IN2 : in std_logic;  Q : out std_logic);
   end component;
   
   component IBUFFX16
      port( INP : in std_logic;  ZN : out std_logic);
   end component;
   
   component DELLN2X2
      port( INP : in std_logic;  Z : out std_logic);
   end component;
   
   component AO22X2
      port( IN1, IN2, IN3, IN4 : in std_logic;  Q : out std_logic);
   end component;
   
   component AND2X4
      port( IN1, IN2 : in std_logic;  Q : out std_logic);
   end component;
   
   component NAND3X4
      port( IN1, IN2, IN3 : in std_logic;  QN : out std_logic);
   end component;
   
   component NAND4X1
      port( IN1, IN2, IN3, IN4 : in std_logic;  QN : out std_logic);
   end component;
   
   component AO221X1
      port( IN1, IN2, IN3, IN4, IN5 : in std_logic;  Q : out std_logic);
   end component;
   
   component OR2X4
      port( IN1, IN2 : in std_logic;  Q : out std_logic);
   end component;
   
   component DELLN1X2
      port( INP : in std_logic;  Z : out std_logic);
   end component;
   
   component AO221X2
      port( IN1, IN2, IN3, IN4, IN5 : in std_logic;  Q : out std_logic);
   end component;
   
   component OR2X2
      port( IN1, IN2 : in std_logic;  Q : out std_logic);
   end component;
   
   component DFFX1
      port( D, CLK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component CryptoCore_1_DW01_cmp6_0
      port( A, B : in std_logic_vector (31 downto 0);  TC : in std_logic;  LT, 
            GT, EQ, LE, GE, NE : out std_logic);
   end component;
   
   component cyclist_ops_RAM_LEN128_DATA_LEN32_1
      port( cyc_state_update_sel, xor_sel, cycd_sel : in std_logic_vector (1 
            downto 0);  extract_sel, addr_sel2 : in std_logic;  ramoutd1 : in 
            std_logic_vector (127 downto 0);  key, bdi_data : in 
            std_logic_vector (31 downto 0);  cu_cd : in std_logic_vector (7 
            downto 0);  dcount_in : in std_logic_vector (1 downto 0);  
            cyc_state_update : out std_logic_vector (127 downto 0);  bdo_out : 
            out std_logic_vector (31 downto 0));
   end component;
   
   component counter_num_bits4_1_1
      port( clk, load, enable : in std_logic;  start_value : in 
            std_logic_vector (3 downto 0);  q : out std_logic_vector (3 downto 
            0));
   end component;
   
   component counter_num_bits5_1
      port( clk, load, enable : in std_logic;  start_value : in 
            std_logic_vector (4 downto 0);  q : out std_logic_vector (4 downto 
            0));
   end component;
   
   component counter_num_bits4_1_0
      port( clk, load, enable : in std_logic;  start_value : in 
            std_logic_vector (3 downto 0);  q : out std_logic_vector (3 downto 
            0));
   end component;
   
   component 
      xoodoo_round_ADDRESS_LEN128_ADDRESS_ENTRIES16_ADDRESS_ENTRIES_BITs4_1
      port( RAMA, RAMB : in std_logic_vector (127 downto 0);  perm_output : out
            std_logic_vector (127 downto 0);  ADDRA, ADDRB : out 
            std_logic_vector (3 downto 0);  RNDCTR : in std_logic_vector (3 
            downto 0);  ins_counter : in std_logic_vector (4 downto 0));
   end component;
   
   component DUAL_PORT_RAM_32_BIT_ADDRESS_LEN128_ADDR_ENTRIES16_ADD_ENT_BITS4_1
      port( RAMADDR1, RAMADDR2 : in std_logic_vector (3 downto 0);  RAMDIN1 : 
            in std_logic_vector (127 downto 0);  RAMDOUT1, RAMDOUT2 : out 
            std_logic_vector (127 downto 0);  RAMWRITE1, clk : in std_logic);
   end component;
   
   component OA21X1
      port( IN1, IN2, IN3 : in std_logic;  Q : out std_logic);
   end component;
   
   component AOI22X1
      port( IN1, IN2, IN3, IN4 : in std_logic;  QN : out std_logic);
   end component;
   
   component AO222X1
      port( IN1, IN2, IN3, IN4, IN5, IN6 : in std_logic;  Q : out std_logic);
   end component;
   
   component OAI21X1
      port( IN1, IN2, IN3 : in std_logic;  QN : out std_logic);
   end component;
   
   component OAI22X1
      port( IN1, IN2, IN3, IN4 : in std_logic;  QN : out std_logic);
   end component;
   
   component OA22X1
      port( IN1, IN2, IN3, IN4 : in std_logic;  Q : out std_logic);
   end component;
   
   component OA222X1
      port( IN1, IN2, IN3, IN4, IN5, IN6 : in std_logic;  Q : out std_logic);
   end component;
   
   signal X_Logic0_port, n265, n266, bdo_29_port, bdo_28_port, bdo_27_port, 
      bdo_26_port, bdo_25_port, bdo_24_port, bdo_23_port, bdo_22_port, 
      bdo_21_port, bdo_20_port, bdo_19_port, bdo_18_port, bdo_17_port, 
      bdo_16_port, bdo_15_port, bdo_14_port, bdo_13_port, bdo_12_port, 
      bdo_11_port, bdo_10_port, bdo_9_port, bdo_8_port, n267, n268, n269, 
      bdo_4_port, n270, bdo_2_port, n271, bdo_0_port, bdo_type_3_port, 
      addrmux2_3_port, addrmux2_2_port, addrmux2_1_port, addrmux2_0_port, 
      perm_addr2_3_port, perm_addr2_2_port, perm_addr2_1_port, 
      perm_addr2_0_port, ramainput_127_port, ramainput_126_port, 
      ramainput_125_port, ramainput_124_port, ramainput_123_port, 
      ramainput_122_port, ramainput_121_port, ramainput_120_port, 
      ramainput_119_port, ramainput_118_port, ramainput_117_port, 
      ramainput_116_port, ramainput_115_port, ramainput_114_port, 
      ramainput_113_port, ramainput_112_port, ramainput_111_port, 
      ramainput_110_port, ramainput_109_port, ramainput_108_port, 
      ramainput_107_port, ramainput_106_port, ramainput_105_port, 
      ramainput_104_port, ramainput_103_port, ramainput_102_port, 
      ramainput_101_port, ramainput_100_port, ramainput_99_port, 
      ramainput_98_port, ramainput_97_port, ramainput_96_port, 
      ramainput_95_port, ramainput_94_port, ramainput_93_port, 
      ramainput_92_port, ramainput_91_port, ramainput_90_port, 
      ramainput_89_port, ramainput_88_port, ramainput_87_port, 
      ramainput_86_port, ramainput_85_port, ramainput_84_port, 
      ramainput_83_port, ramainput_82_port, ramainput_81_port, 
      ramainput_80_port, ramainput_79_port, ramainput_78_port, 
      ramainput_77_port, ramainput_76_port, ramainput_75_port, 
      ramainput_74_port, ramainput_73_port, ramainput_72_port, 
      ramainput_71_port, ramainput_70_port, ramainput_69_port, 
      ramainput_68_port, ramainput_67_port, ramainput_66_port, 
      ramainput_65_port, ramainput_64_port, ramainput_63_port, 
      ramainput_62_port, ramainput_61_port, ramainput_60_port, 
      ramainput_59_port, ramainput_58_port, ramainput_57_port, 
      ramainput_56_port, ramainput_55_port, ramainput_54_port, 
      ramainput_53_port, ramainput_52_port, ramainput_51_port, 
      ramainput_50_port, ramainput_49_port, ramainput_48_port, 
      ramainput_47_port, ramainput_46_port, ramainput_45_port, 
      ramainput_44_port, ramainput_43_port, ramainput_42_port, 
      ramainput_41_port, ramainput_40_port, ramainput_39_port, 
      ramainput_38_port, ramainput_37_port, ramainput_36_port, 
      ramainput_35_port, ramainput_34_port, ramainput_33_port, 
      ramainput_32_port, ramainput_31_port, ramainput_30_port, 
      ramainput_29_port, ramainput_28_port, ramainput_27_port, 
      ramainput_26_port, ramainput_25_port, ramainput_24_port, 
      ramainput_23_port, ramainput_22_port, ramainput_21_port, 
      ramainput_20_port, ramainput_19_port, ramainput_18_port, 
      ramainput_17_port, ramainput_16_port, ramainput_15_port, 
      ramainput_14_port, ramainput_13_port, ramainput_12_port, 
      ramainput_11_port, ramainput_10_port, ramainput_9_port, ramainput_8_port,
      ramainput_7_port, ramainput_6_port, ramainput_5_port, ramainput_4_port, 
      ramainput_3_port, ramainput_2_port, ramainput_1_port, ramainput_0_port, 
      ramout1_127_port, ramout1_126_port, ramout1_125_port, ramout1_124_port, 
      ramout1_123_port, ramout1_122_port, ramout1_121_port, ramout1_120_port, 
      ramout1_119_port, ramout1_118_port, ramout1_117_port, ramout1_116_port, 
      ramout1_115_port, ramout1_114_port, ramout1_113_port, ramout1_112_port, 
      ramout1_111_port, ramout1_110_port, ramout1_109_port, ramout1_108_port, 
      ramout1_107_port, ramout1_106_port, ramout1_105_port, ramout1_104_port, 
      ramout1_103_port, ramout1_102_port, ramout1_101_port, ramout1_100_port, 
      ramout1_99_port, ramout1_98_port, ramout1_97_port, ramout1_96_port, 
      ramout1_95_port, ramout1_94_port, ramout1_93_port, ramout1_92_port, 
      ramout1_91_port, ramout1_90_port, ramout1_89_port, ramout1_88_port, 
      ramout1_87_port, ramout1_86_port, ramout1_85_port, ramout1_84_port, 
      ramout1_83_port, ramout1_82_port, ramout1_81_port, ramout1_80_port, 
      ramout1_79_port, ramout1_78_port, ramout1_77_port, ramout1_76_port, 
      ramout1_75_port, ramout1_74_port, ramout1_73_port, ramout1_72_port, 
      ramout1_71_port, ramout1_70_port, ramout1_69_port, ramout1_68_port, 
      ramout1_67_port, ramout1_66_port, ramout1_65_port, ramout1_64_port, 
      ramout1_63_port, ramout1_62_port, ramout1_61_port, ramout1_60_port, 
      ramout1_59_port, ramout1_58_port, ramout1_57_port, ramout1_56_port, 
      ramout1_55_port, ramout1_54_port, ramout1_53_port, ramout1_52_port, 
      ramout1_51_port, ramout1_50_port, ramout1_49_port, ramout1_48_port, 
      ramout1_47_port, ramout1_46_port, ramout1_45_port, ramout1_44_port, 
      ramout1_43_port, ramout1_42_port, ramout1_41_port, ramout1_40_port, 
      ramout1_39_port, ramout1_38_port, ramout1_37_port, ramout1_36_port, 
      ramout1_35_port, ramout1_34_port, ramout1_33_port, ramout1_32_port, 
      ramout1_31_port, ramout1_30_port, ramout1_29_port, ramout1_28_port, 
      ramout1_27_port, ramout1_26_port, ramout1_25_port, ramout1_24_port, 
      ramout1_23_port, ramout1_22_port, ramout1_21_port, ramout1_20_port, 
      ramout1_19_port, ramout1_18_port, ramout1_17_port, ramout1_16_port, 
      ramout1_15_port, ramout1_14_port, ramout1_13_port, ramout1_12_port, 
      ramout1_11_port, ramout1_10_port, ramout1_9_port, ramout1_8_port, 
      ramout1_7_port, ramout1_6_port, ramout1_5_port, ramout1_4_port, 
      ramout1_3_port, ramout1_2_port, ramout1_1_port, ramout1_0_port, 
      ramout2_127_port, ramout2_126_port, ramout2_125_port, ramout2_124_port, 
      ramout2_123_port, ramout2_122_port, ramout2_121_port, ramout2_120_port, 
      ramout2_119_port, ramout2_118_port, ramout2_117_port, ramout2_116_port, 
      ramout2_115_port, ramout2_114_port, ramout2_113_port, ramout2_112_port, 
      ramout2_111_port, ramout2_110_port, ramout2_109_port, ramout2_108_port, 
      ramout2_107_port, ramout2_106_port, ramout2_105_port, ramout2_104_port, 
      ramout2_103_port, ramout2_102_port, ramout2_101_port, ramout2_100_port, 
      ramout2_99_port, ramout2_98_port, ramout2_97_port, ramout2_96_port, 
      ramout2_95_port, ramout2_94_port, ramout2_93_port, ramout2_92_port, 
      ramout2_91_port, ramout2_90_port, ramout2_89_port, ramout2_88_port, 
      ramout2_87_port, ramout2_86_port, ramout2_85_port, ramout2_84_port, 
      ramout2_83_port, ramout2_82_port, ramout2_81_port, ramout2_80_port, 
      ramout2_79_port, ramout2_78_port, ramout2_77_port, ramout2_76_port, 
      ramout2_75_port, ramout2_74_port, ramout2_73_port, ramout2_72_port, 
      ramout2_71_port, ramout2_70_port, ramout2_69_port, ramout2_68_port, 
      ramout2_67_port, ramout2_66_port, ramout2_65_port, ramout2_64_port, 
      ramout2_63_port, ramout2_62_port, ramout2_61_port, ramout2_60_port, 
      ramout2_59_port, ramout2_58_port, ramout2_57_port, ramout2_56_port, 
      ramout2_55_port, ramout2_54_port, ramout2_53_port, ramout2_52_port, 
      ramout2_51_port, ramout2_50_port, ramout2_49_port, ramout2_48_port, 
      ramout2_47_port, ramout2_46_port, ramout2_45_port, ramout2_44_port, 
      ramout2_43_port, ramout2_42_port, ramout2_41_port, ramout2_40_port, 
      ramout2_39_port, ramout2_38_port, ramout2_37_port, ramout2_36_port, 
      ramout2_35_port, ramout2_34_port, ramout2_33_port, ramout2_32_port, 
      ramout2_31_port, ramout2_30_port, ramout2_29_port, ramout2_28_port, 
      ramout2_27_port, ramout2_26_port, ramout2_25_port, ramout2_24_port, 
      ramout2_23_port, ramout2_22_port, ramout2_21_port, ramout2_20_port, 
      ramout2_19_port, ramout2_18_port, ramout2_17_port, ramout2_16_port, 
      ramout2_15_port, ramout2_14_port, ramout2_13_port, ramout2_12_port, 
      ramout2_11_port, ramout2_10_port, ramout2_9_port, ramout2_8_port, 
      ramout2_7_port, ramout2_6_port, ramout2_5_port, ramout2_4_port, 
      ramout2_3_port, ramout2_2_port, ramout2_1_port, ramout2_0_port, ramwrite,
      perm_output_127_port, perm_output_126_port, perm_output_125_port, 
      perm_output_124_port, perm_output_123_port, perm_output_122_port, 
      perm_output_121_port, perm_output_120_port, perm_output_119_port, 
      perm_output_118_port, perm_output_117_port, perm_output_116_port, 
      perm_output_115_port, perm_output_114_port, perm_output_113_port, 
      perm_output_112_port, perm_output_111_port, perm_output_110_port, 
      perm_output_109_port, perm_output_108_port, perm_output_107_port, 
      perm_output_106_port, perm_output_105_port, perm_output_104_port, 
      perm_output_103_port, perm_output_102_port, perm_output_101_port, 
      perm_output_100_port, perm_output_99_port, perm_output_98_port, 
      perm_output_97_port, perm_output_96_port, perm_output_95_port, 
      perm_output_94_port, perm_output_93_port, perm_output_92_port, 
      perm_output_91_port, perm_output_90_port, perm_output_89_port, 
      perm_output_88_port, perm_output_87_port, perm_output_86_port, 
      perm_output_85_port, perm_output_84_port, perm_output_83_port, 
      perm_output_82_port, perm_output_81_port, perm_output_80_port, 
      perm_output_79_port, perm_output_78_port, perm_output_77_port, 
      perm_output_76_port, perm_output_75_port, perm_output_74_port, 
      perm_output_73_port, perm_output_72_port, perm_output_71_port, 
      perm_output_70_port, perm_output_69_port, perm_output_68_port, 
      perm_output_67_port, perm_output_66_port, perm_output_65_port, 
      perm_output_64_port, perm_output_63_port, perm_output_62_port, 
      perm_output_61_port, perm_output_60_port, perm_output_59_port, 
      perm_output_58_port, perm_output_57_port, perm_output_56_port, 
      perm_output_55_port, perm_output_54_port, perm_output_53_port, 
      perm_output_52_port, perm_output_51_port, perm_output_50_port, 
      perm_output_49_port, perm_output_48_port, perm_output_47_port, 
      perm_output_46_port, perm_output_45_port, perm_output_44_port, 
      perm_output_43_port, perm_output_42_port, perm_output_41_port, 
      perm_output_40_port, perm_output_39_port, perm_output_38_port, 
      perm_output_37_port, perm_output_36_port, perm_output_35_port, 
      perm_output_34_port, perm_output_33_port, perm_output_32_port, 
      perm_output_31_port, perm_output_30_port, perm_output_29_port, 
      perm_output_28_port, perm_output_27_port, perm_output_26_port, 
      perm_output_25_port, perm_output_24_port, perm_output_23_port, 
      perm_output_22_port, perm_output_21_port, perm_output_20_port, 
      perm_output_19_port, perm_output_18_port, perm_output_17_port, 
      perm_output_16_port, perm_output_15_port, perm_output_14_port, 
      perm_output_13_port, perm_output_12_port, perm_output_11_port, 
      perm_output_10_port, perm_output_9_port, perm_output_8_port, 
      perm_output_7_port, perm_output_6_port, perm_output_5_port, 
      perm_output_4_port, perm_output_3_port, perm_output_2_port, 
      perm_output_1_port, perm_output_0_port, cyc_state_update_127_port, 
      cyc_state_update_126_port, cyc_state_update_125_port, 
      cyc_state_update_124_port, cyc_state_update_123_port, 
      cyc_state_update_122_port, cyc_state_update_121_port, 
      cyc_state_update_120_port, cyc_state_update_119_port, 
      cyc_state_update_118_port, cyc_state_update_117_port, 
      cyc_state_update_116_port, cyc_state_update_115_port, 
      cyc_state_update_114_port, cyc_state_update_113_port, 
      cyc_state_update_112_port, cyc_state_update_111_port, 
      cyc_state_update_110_port, cyc_state_update_109_port, 
      cyc_state_update_108_port, cyc_state_update_107_port, 
      cyc_state_update_106_port, cyc_state_update_105_port, 
      cyc_state_update_104_port, cyc_state_update_103_port, 
      cyc_state_update_102_port, cyc_state_update_101_port, 
      cyc_state_update_100_port, cyc_state_update_99_port, 
      cyc_state_update_98_port, cyc_state_update_97_port, 
      cyc_state_update_96_port, cyc_state_update_95_port, 
      cyc_state_update_94_port, cyc_state_update_93_port, 
      cyc_state_update_92_port, cyc_state_update_91_port, 
      cyc_state_update_90_port, cyc_state_update_89_port, 
      cyc_state_update_88_port, cyc_state_update_87_port, 
      cyc_state_update_86_port, cyc_state_update_85_port, 
      cyc_state_update_84_port, cyc_state_update_83_port, 
      cyc_state_update_82_port, cyc_state_update_81_port, 
      cyc_state_update_80_port, cyc_state_update_79_port, 
      cyc_state_update_78_port, cyc_state_update_77_port, 
      cyc_state_update_76_port, cyc_state_update_75_port, 
      cyc_state_update_74_port, cyc_state_update_73_port, 
      cyc_state_update_72_port, cyc_state_update_71_port, 
      cyc_state_update_70_port, cyc_state_update_69_port, 
      cyc_state_update_68_port, cyc_state_update_67_port, 
      cyc_state_update_66_port, cyc_state_update_65_port, 
      cyc_state_update_64_port, cyc_state_update_63_port, 
      cyc_state_update_62_port, cyc_state_update_61_port, 
      cyc_state_update_60_port, cyc_state_update_59_port, 
      cyc_state_update_58_port, cyc_state_update_57_port, 
      cyc_state_update_56_port, cyc_state_update_55_port, 
      cyc_state_update_54_port, cyc_state_update_53_port, 
      cyc_state_update_52_port, cyc_state_update_51_port, 
      cyc_state_update_50_port, cyc_state_update_49_port, 
      cyc_state_update_48_port, cyc_state_update_47_port, 
      cyc_state_update_46_port, cyc_state_update_45_port, 
      cyc_state_update_44_port, cyc_state_update_43_port, 
      cyc_state_update_42_port, cyc_state_update_41_port, 
      cyc_state_update_40_port, cyc_state_update_39_port, 
      cyc_state_update_38_port, cyc_state_update_37_port, 
      cyc_state_update_36_port, cyc_state_update_35_port, 
      cyc_state_update_34_port, cyc_state_update_33_port, 
      cyc_state_update_32_port, cyc_state_update_31_port, 
      cyc_state_update_30_port, cyc_state_update_29_port, 
      cyc_state_update_28_port, cyc_state_update_27_port, 
      cyc_state_update_26_port, cyc_state_update_25_port, 
      cyc_state_update_24_port, cyc_state_update_23_port, 
      cyc_state_update_22_port, cyc_state_update_21_port, 
      cyc_state_update_20_port, cyc_state_update_19_port, 
      cyc_state_update_18_port, cyc_state_update_17_port, 
      cyc_state_update_16_port, cyc_state_update_15_port, 
      cyc_state_update_14_port, cyc_state_update_13_port, 
      cyc_state_update_12_port, cyc_state_update_11_port, 
      cyc_state_update_10_port, cyc_state_update_9_port, 
      cyc_state_update_8_port, cyc_state_update_7_port, cyc_state_update_6_port
      , cyc_state_update_5_port, cyc_state_update_4_port, 
      cyc_state_update_3_port, cyc_state_update_2_port, cyc_state_update_1_port
      , cyc_state_update_0_port, addr_sel_1_port, perm_addr_3_port, 
      perm_addr_2_port, perm_addr_1_port, perm_addr_0_port, dcount_3_port, 
      dcount_2_port, dcount_1_port, dcount_0_port, rnd_counter_3_port, 
      rnd_counter_2_port, rnd_counter_1_port, rnd_counter_0_port, 
      ins_counter_4_port, ins_counter_3_port, ins_counter_2_port, 
      ins_counter_1_port, ins_counter_0_port, load_rnd, en_rnd, load_ins, 
      en_ins, ins_start_value_4_port, ins_start_value_3_port, ins_start_value_0
      , load_dcount, en_dcount, dcount_start_value_3, 
      cyc_state_update_sel_1_port, cyc_state_update_sel_0_port, xor_sel_1_port,
      cycd_sel_1_port, cycd_sel_0_port, extract_sel, cu_cd_s_6_port, cu_cd_s_1,
      calling_state_2_port, calling_state_1_port, calling_state_0_port, N72, 
      N73, cyc_s_2_port, cyc_s_1_port, cyc_s_0_port, key_update_internal_0_port
      , decrypt_op_s, gtr_one_perm, N103, N275, tag_verified, N305, N306, N307,
      n1, n31, n44, n45, n46, n51, n52, n53, n54, n64, n65, n66, n67, n68, n69,
      n70, n71, n72_port, n73_port, n74, n75, n76, n77, n78, n79, n80, n81, n82
      , n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, 
      n97, n98, n99, n100, n101, n102, n103_port, n104, n105, n106, n107, n108,
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195, n196, n198, n199, n204, n205, n206, n207, n208, n209, 
      n210, n211, n212, n213, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, 
      n13, n14, n15, n16, n17, n18, n19, n20, n21, bdo_3_port, bdo_1_port, 
      bdo_30_port, bdo_5_port, n26, bdo_7_port, bdo_6_port, n29, n30, n32, n33,
      n34, n35, n36, n37, key_ready_port, n39, n40, n41, n42, bdo_31_port, n47,
      n48, n49, n50, n55, n56, n57, n58, n59, n60, n61, n62, n63, n197, n200, 
      n201, n202, n203, n214, n215, n216, n217, n218, n219, n220, n221, n222, 
      n223, n224, n225, n226, n227, bdo_type_0_port, n229, n230, n231, n232, 
      n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, 
      n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, 
      n257, n258, n259, n260, n261, n262, n263, n264, n_3222, n_3223, n_3224, 
      n_3225, n_3226, n_3227, n_3228, n_3229, n_3230 : std_logic;

begin
   key_ready <= key_ready_port;
   bdo <= ( bdo_31_port, bdo_30_port, bdo_29_port, bdo_28_port, bdo_27_port, 
      bdo_26_port, bdo_25_port, bdo_24_port, bdo_23_port, bdo_22_port, 
      bdo_21_port, bdo_20_port, bdo_19_port, bdo_18_port, bdo_17_port, 
      bdo_16_port, bdo_15_port, bdo_14_port, bdo_13_port, bdo_12_port, 
      bdo_11_port, bdo_10_port, bdo_9_port, bdo_8_port, bdo_7_port, bdo_6_port,
      bdo_5_port, bdo_4_port, bdo_3_port, bdo_2_port, bdo_1_port, bdo_0_port );
   bdo_type <= ( bdo_type_3_port, extract_sel, X_Logic0_port, bdo_type_0_port )
      ;
   
   X_Logic0_port <= '0';
   n1 <= '0';
   decrypt_op_s_reg : DFFX1 port map( D => n213, CLK => n40, Q => decrypt_op_s,
                           QN => n54);
   key_update_internal_reg_1_inst : DFFX1 port map( D => n211, CLK => n40, Q =>
                           n33, QN => n31);
   calling_state_reg_2_inst : DFFX1 port map( D => n207, CLK => n40, Q => 
                           calling_state_2_port, QN => n51);
   calling_state_reg_1_inst : DFFX1 port map( D => n206, CLK => n40, Q => 
                           calling_state_1_port, QN => n52);
   cyc_s_reg_0_inst : DFFX1 port map( D => n210, CLK => n40, Q => cyc_s_0_port,
                           QN => n46);
   calling_state_reg_0_inst : DFFX1 port map( D => n205, CLK => n40, Q => 
                           calling_state_0_port, QN => n_3222);
   gtr_one_perm_reg : DFFX1 port map( D => n204, CLK => n40, Q => gtr_one_perm,
                           QN => n53);
   msg_auth_valid_reg : DFFX1 port map( D => N306, CLK => n40, Q => 
                           msg_auth_valid, QN => n_3223);
   key_update_internal_reg_0_inst : DFFX1 port map( D => n208, CLK => n40, Q =>
                           key_update_internal_0_port, QN => n34);
   tag_verified_reg : DFFX1 port map( D => N307, CLK => n40, Q => tag_verified,
                           QN => n_3224);
   msg_auth_reg : DFFX1 port map( D => N305, CLK => n40, Q => msg_auth, QN => 
                           n_3225);
   U123 : NAND4X0 port map( IN1 => n257, IN2 => n65, IN3 => n66, IN4 => n67, QN
                           => ramwrite);
   U124 : OA21X1 port map( IN1 => n238, IN2 => n68, IN3 => n69, Q => n67);
   U177 : AO22X1 port map( IN1 => perm_output_52_port, IN2 => n220, IN3 => 
                           cyc_state_update_52_port, IN4 => n55, Q => 
                           ramainput_52_port);
   U194 : AO22X1 port map( IN1 => perm_output_37_port, IN2 => n215, IN3 => 
                           cyc_state_update_37_port, IN4 => n56, Q => 
                           ramainput_37_port);
   U255 : AO22X1 port map( IN1 => calling_state_0_port, IN2 => n76, IN3 => n77,
                           IN4 => n72_port, Q => n205);
   U257 : OAI21X1 port map( IN1 => n76, IN2 => n72_port, IN3 => 
                           calling_state_1_port, QN => n78);
   U258 : NAND3X0 port map( IN1 => n83, IN2 => n264, IN3 => n84, QN => n82);
   U260 : OA21X1 port map( IN1 => n86, IN2 => n87, IN3 => n264, Q => n85);
   U261 : NAND4X0 port map( IN1 => n75, IN2 => n89, IN3 => n90, IN4 => n246, QN
                           => n88);
   U262 : AO22X1 port map( IN1 => key_update_internal_0_port, IN2 => n92, IN3 
                           => n93, IN4 => key_update, Q => n208);
   U263 : NAND3X0 port map( IN1 => n95, IN2 => n96, IN3 => n248, QN => n92);
   U264 : AO22X1 port map( IN1 => n98, IN2 => cyc_s_1_port, IN3 => n99, IN4 => 
                           n100, Q => n209);
   U265 : NAND3X0 port map( IN1 => n9, IN2 => n102, IN3 => n103_port, QN => 
                           n100);
   U266 : OA22X1 port map( IN1 => n104, IN2 => n105, IN3 => n41, IN4 => n83, Q 
                           => n103_port);
   U267 : AO22X1 port map( IN1 => n98, IN2 => cyc_s_0_port, IN3 => n99, IN4 => 
                           n106, Q => n210);
   U268 : NAND4X0 port map( IN1 => n107, IN2 => n81, IN3 => n108, IN4 => n109, 
                           QN => n106);
   U269 : OA222X1 port map( IN1 => n110, IN2 => n111, IN3 => n112, IN4 => n46, 
                           IN5 => n105, IN6 => n258, Q => n109);
   U270 : OA21X1 port map( IN1 => n231, IN2 => n244, IN3 => n102, Q => n112);
   U271 : AND3X1 port map( IN1 => n113, IN2 => n68, IN3 => n114, Q => n102);
   U272 : OA22X1 port map( IN1 => n259, IN2 => n116, IN3 => n117, IN4 => n118, 
                           Q => n110);
   U273 : AND3X1 port map( IN1 => n119, IN2 => n120, IN3 => n121, Q => n117);
   U274 : NAND4X0 port map( IN1 => dcount_3_port, IN2 => dcount_1_port, IN3 => 
                           n122, IN4 => bdi_valid, QN => n120);
   U275 : AND3X1 port map( IN1 => n123, IN2 => n124, IN3 => n125, Q => n116);
   U276 : NAND3X0 port map( IN1 => dcount_0_port, IN2 => n126, IN3 => n127, QN 
                           => n125);
   U277 : NAND3X0 port map( IN1 => n233, IN2 => n250, IN3 => n129, QN => n107);
   U278 : OAI21X1 port map( IN1 => n130, IN2 => n31, IN3 => n131, QN => n211);
   U280 : OA21X1 port map( IN1 => n86, IN2 => n41, IN3 => n248, Q => n130);
   U282 : NOR3X0 port map( IN1 => n250, IN2 => n8, IN3 => n133, QN => n75);
   U283 : AO22X1 port map( IN1 => n98, IN2 => cyc_s_2_port, IN3 => n99, IN4 => 
                           n134, Q => n212);
   U284 : NAND4X0 port map( IN1 => n114, IN2 => n135, IN3 => n9, IN4 => n136, 
                           QN => n134);
   U285 : NOR3X0 port map( IN1 => n254, IN2 => n128, IN3 => n8, QN => n136);
   U286 : AOI22X1 port map( IN1 => n249, IN2 => n138, IN3 => n139, IN4 => n140,
                           QN => n114);
   U287 : OR2X1 port map( IN1 => bdo_type_3_port, IN2 => n141, Q => n139);
   U288 : AOI21X1 port map( IN1 => n143, IN2 => n246, IN3 => rst, QN => n98);
   U289 : AO22X1 port map( IN1 => cyc_s_0_port, IN2 => n144, IN3 => n145, IN4 
                           => n46, Q => n143);
   U290 : NAND3X0 port map( IN1 => n148, IN2 => n149, IN3 => decrypt_op_s, QN 
                           => n144);
   U291 : OAI22X1 port map( IN1 => n54, IN2 => n150, IN3 => rst, IN4 => n151, 
                           QN => n213);
   U292 : OA21X1 port map( IN1 => n152, IN2 => n54, IN3 => n153, Q => n151);
   U293 : NAND3X0 port map( IN1 => n152, IN2 => n150, IN3 => decrypt_in, QN => 
                           n153);
   U296 : NAND4X0 port map( IN1 => n91, IN2 => n3, IN3 => n90, IN4 => n236, QN 
                           => load_ins);
   U297 : NAND4X0 port map( IN1 => n158, IN2 => n160, IN3 => n161, IN4 => n156,
                           QN => load_dcount);
   U300 : OR2X1 port map( IN1 => n236, IN2 => n115, Q => n105);
   U301 : OR2X1 port map( IN1 => ins_start_value_0, IN2 => 
                           ins_start_value_3_port, Q => ins_start_value_4_port)
                           ;
   U302 : NOR3X0 port map( IN1 => n146, IN2 => key_update, IN3 => n90, QN => 
                           ins_start_value_3_port);
   U303 : NAND4X0 port map( IN1 => rnd_counter_3_port, IN2 => 
                           rnd_counter_1_port, IN3 => rnd_counter_0_port, IN4 
                           => n237, QN => n115);
   U304 : NOR3X0 port map( IN1 => calling_state_0_port, IN2 => 
                           calling_state_1_port, IN3 => n51, QN => n104);
   U305 : NOR3X0 port map( IN1 => n165, IN2 => bdo_type_3_port, IN3 => n166, QN
                           => n164);
   U306 : NAND3X0 port map( IN1 => ins_counter_4_port, IN2 => 
                           ins_counter_2_port, IN3 => n169, QN => n138);
   U307 : NOR3X0 port map( IN1 => ins_counter_0_port, IN2 => ins_counter_3_port
                           , IN3 => ins_counter_1_port, QN => n169);
   U308 : NAND4X0 port map( IN1 => n170, IN2 => n171, IN3 => n172, IN4 => n173,
                           QN => en_dcount);
   U309 : NAND3X0 port map( IN1 => n173, IN2 => n91, IN3 => n174, QN => 
                           dcount_start_value_3);
   U310 : NAND4X0 port map( IN1 => n175, IN2 => n234, IN3 => dcount_1_port, IN4
                           => n176, QN => n97);
   U312 : NAND4X0 port map( IN1 => n127, IN2 => key_ready_port, IN3 => n175, 
                           IN4 => n232, QN => n179);
   U313 : NOR3X0 port map( IN1 => dcount_1_port, IN2 => dcount_3_port, IN3 => 
                           n234, QN => n127);
   U314 : OAI21X1 port map( IN1 => n175, IN2 => n246, IN3 => n178, QN => 
                           cyc_state_update_sel_0_port);
   U315 : NAND4X0 port map( IN1 => n254, IN2 => n52, IN3 => n51, IN4 => n53, QN
                           => n65);
   U316 : NAND4X0 port map( IN1 => n180, IN2 => n256, IN3 => 
                           calling_state_1_port, IN4 => n53, QN => n66);
   U317 : NOR3X0 port map( IN1 => n137, IN2 => gtr_one_perm, IN3 => n156, QN =>
                           cu_cd_s_6_port);
   U318 : AO21X1 port map( IN1 => bdi_valid_bytes(3), IN2 => extract_sel, IN3 
                           => bdo_type_3_port, Q => bdo_valid_bytes(3));
   U319 : AO21X1 port map( IN1 => bdi_valid_bytes(2), IN2 => extract_sel, IN3 
                           => bdo_type_3_port, Q => bdo_valid_bytes(2));
   U320 : AO21X1 port map( IN1 => bdi_valid_bytes(1), IN2 => extract_sel, IN3 
                           => bdo_type_3_port, Q => bdo_valid_bytes(1));
   U321 : AO21X1 port map( IN1 => bdi_valid_bytes(0), IN2 => extract_sel, IN3 
                           => bdo_type_3_port, Q => bdo_valid_bytes(0));
   U323 : AO21X1 port map( IN1 => n230, IN2 => n184, IN3 => n165, Q => n183);
   U324 : AO21X1 port map( IN1 => n182, IN2 => n36, IN3 => n165, Q => 
                           extract_sel);
   U326 : AND2X1 port map( IN1 => n186, IN2 => n184, Q => n182);
   U328 : AO222X1 port map( IN1 => n189, IN2 => n184, IN3 => n190, IN4 => 
                           bdi_type(3), IN5 => bdi_type(0), IN6 => n191, Q => 
                           n73_port);
   U329 : OA21X1 port map( IN1 => n192, IN2 => n193, IN3 => n263, Q => n190);
   U330 : AND3X1 port map( IN1 => bdi_type(0), IN2 => n185, IN3 => bdi_type(2),
                           Q => n193);
   U331 : NOR3X0 port map( IN1 => n137, IN2 => bdi_type(2), IN3 => bdi_type(0),
                           QN => n192);
   U333 : AO22X1 port map( IN1 => N72, IN2 => n259, IN3 => N73, IN4 => 
                           calling_state_1_port, Q => n187);
   U334 : AOI22X1 port map( IN1 => n250, IN2 => n70, IN3 => n243, IN4 => n141, 
                           QN => n170);
   U335 : AO221X1 port map( IN1 => n191, IN2 => n194, IN3 => n181, IN4 => n118,
                           IN5 => n129, Q => n70);
   U337 : AND2X1 port map( IN1 => n195, IN2 => n123, Q => n181);
   U338 : AO21X1 port map( IN1 => n119, IN2 => n261, IN3 => n184, Q => n123);
   U339 : NOR3X0 port map( IN1 => bdi_type(1), IN2 => bdi_type(3), IN3 => n262,
                           QN => n184);
   U340 : AO22X1 port map( IN1 => n196, IN2 => bdo_ready, IN3 => n126, IN4 => 
                           n124, Q => n195);
   U341 : AND2X1 port map( IN1 => bdo_ready, IN2 => bdi_valid, Q => n126);
   U342 : AO21X1 port map( IN1 => n121, IN2 => bdi_valid, IN3 => n196, Q => 
                           n194);
   U343 : AND4X1 port map( IN1 => bdi_size(2), IN2 => bdi_eot, IN3 => n188, IN4
                           => bdi_valid, Q => n196);
   U344 : AND2X1 port map( IN1 => n119, IN2 => n259, Q => n191);
   U346 : NOR3X0 port map( IN1 => bdi_type(2), IN2 => bdi_type(3), IN3 => 
                           bdi_type(1), QN => n119);
   U353 : OA21X1 port map( IN1 => n74, IN2 => n32, IN3 => n156, Q => n101);
   U358 : AND3X1 port map( IN1 => n173, IN2 => n41, IN3 => n142, Q => n69);
   U362 : AND3X1 port map( IN1 => N306, IN2 => n229, IN3 => tag_verified, Q => 
                           N305);
   U363 : AND4X1 port map( IN1 => n243, IN2 => n141, IN3 => n233, IN4 => n264, 
                           Q => N306);
   U364 : AND3X1 port map( IN1 => n234, IN2 => n235, IN3 => dcount_1_port, Q =>
                           n163);
   UUT_RAM : DUAL_PORT_RAM_32_BIT_ADDRESS_LEN128_ADDR_ENTRIES16_ADD_ENT_BITS4_1
                           port map( RAMADDR1(3) => addrmux2_3_port, 
                           RAMADDR1(2) => addrmux2_2_port, RAMADDR1(1) => 
                           addrmux2_1_port, RAMADDR1(0) => addrmux2_0_port, 
                           RAMADDR2(3) => perm_addr2_3_port, RAMADDR2(2) => 
                           perm_addr2_2_port, RAMADDR2(1) => perm_addr2_1_port,
                           RAMADDR2(0) => perm_addr2_0_port, RAMDIN1(127) => 
                           ramainput_127_port, RAMDIN1(126) => 
                           ramainput_126_port, RAMDIN1(125) => 
                           ramainput_125_port, RAMDIN1(124) => 
                           ramainput_124_port, RAMDIN1(123) => 
                           ramainput_123_port, RAMDIN1(122) => 
                           ramainput_122_port, RAMDIN1(121) => 
                           ramainput_121_port, RAMDIN1(120) => 
                           ramainput_120_port, RAMDIN1(119) => 
                           ramainput_119_port, RAMDIN1(118) => 
                           ramainput_118_port, RAMDIN1(117) => 
                           ramainput_117_port, RAMDIN1(116) => 
                           ramainput_116_port, RAMDIN1(115) => 
                           ramainput_115_port, RAMDIN1(114) => 
                           ramainput_114_port, RAMDIN1(113) => 
                           ramainput_113_port, RAMDIN1(112) => 
                           ramainput_112_port, RAMDIN1(111) => 
                           ramainput_111_port, RAMDIN1(110) => 
                           ramainput_110_port, RAMDIN1(109) => 
                           ramainput_109_port, RAMDIN1(108) => 
                           ramainput_108_port, RAMDIN1(107) => 
                           ramainput_107_port, RAMDIN1(106) => 
                           ramainput_106_port, RAMDIN1(105) => 
                           ramainput_105_port, RAMDIN1(104) => 
                           ramainput_104_port, RAMDIN1(103) => 
                           ramainput_103_port, RAMDIN1(102) => 
                           ramainput_102_port, RAMDIN1(101) => 
                           ramainput_101_port, RAMDIN1(100) => 
                           ramainput_100_port, RAMDIN1(99) => ramainput_99_port
                           , RAMDIN1(98) => ramainput_98_port, RAMDIN1(97) => 
                           ramainput_97_port, RAMDIN1(96) => ramainput_96_port,
                           RAMDIN1(95) => ramainput_95_port, RAMDIN1(94) => 
                           ramainput_94_port, RAMDIN1(93) => ramainput_93_port,
                           RAMDIN1(92) => ramainput_92_port, RAMDIN1(91) => 
                           ramainput_91_port, RAMDIN1(90) => ramainput_90_port,
                           RAMDIN1(89) => ramainput_89_port, RAMDIN1(88) => 
                           ramainput_88_port, RAMDIN1(87) => ramainput_87_port,
                           RAMDIN1(86) => ramainput_86_port, RAMDIN1(85) => 
                           ramainput_85_port, RAMDIN1(84) => ramainput_84_port,
                           RAMDIN1(83) => ramainput_83_port, RAMDIN1(82) => 
                           ramainput_82_port, RAMDIN1(81) => ramainput_81_port,
                           RAMDIN1(80) => ramainput_80_port, RAMDIN1(79) => 
                           ramainput_79_port, RAMDIN1(78) => ramainput_78_port,
                           RAMDIN1(77) => ramainput_77_port, RAMDIN1(76) => 
                           ramainput_76_port, RAMDIN1(75) => ramainput_75_port,
                           RAMDIN1(74) => ramainput_74_port, RAMDIN1(73) => 
                           ramainput_73_port, RAMDIN1(72) => ramainput_72_port,
                           RAMDIN1(71) => ramainput_71_port, RAMDIN1(70) => 
                           ramainput_70_port, RAMDIN1(69) => ramainput_69_port,
                           RAMDIN1(68) => ramainput_68_port, RAMDIN1(67) => 
                           ramainput_67_port, RAMDIN1(66) => ramainput_66_port,
                           RAMDIN1(65) => ramainput_65_port, RAMDIN1(64) => 
                           ramainput_64_port, RAMDIN1(63) => ramainput_63_port,
                           RAMDIN1(62) => ramainput_62_port, RAMDIN1(61) => 
                           ramainput_61_port, RAMDIN1(60) => ramainput_60_port,
                           RAMDIN1(59) => ramainput_59_port, RAMDIN1(58) => 
                           ramainput_58_port, RAMDIN1(57) => ramainput_57_port,
                           RAMDIN1(56) => ramainput_56_port, RAMDIN1(55) => 
                           ramainput_55_port, RAMDIN1(54) => ramainput_54_port,
                           RAMDIN1(53) => ramainput_53_port, RAMDIN1(52) => 
                           ramainput_52_port, RAMDIN1(51) => ramainput_51_port,
                           RAMDIN1(50) => ramainput_50_port, RAMDIN1(49) => 
                           ramainput_49_port, RAMDIN1(48) => ramainput_48_port,
                           RAMDIN1(47) => ramainput_47_port, RAMDIN1(46) => 
                           ramainput_46_port, RAMDIN1(45) => ramainput_45_port,
                           RAMDIN1(44) => ramainput_44_port, RAMDIN1(43) => 
                           ramainput_43_port, RAMDIN1(42) => ramainput_42_port,
                           RAMDIN1(41) => ramainput_41_port, RAMDIN1(40) => 
                           ramainput_40_port, RAMDIN1(39) => ramainput_39_port,
                           RAMDIN1(38) => ramainput_38_port, RAMDIN1(37) => 
                           ramainput_37_port, RAMDIN1(36) => ramainput_36_port,
                           RAMDIN1(35) => ramainput_35_port, RAMDIN1(34) => 
                           ramainput_34_port, RAMDIN1(33) => ramainput_33_port,
                           RAMDIN1(32) => ramainput_32_port, RAMDIN1(31) => 
                           ramainput_31_port, RAMDIN1(30) => ramainput_30_port,
                           RAMDIN1(29) => ramainput_29_port, RAMDIN1(28) => 
                           ramainput_28_port, RAMDIN1(27) => ramainput_27_port,
                           RAMDIN1(26) => ramainput_26_port, RAMDIN1(25) => 
                           ramainput_25_port, RAMDIN1(24) => ramainput_24_port,
                           RAMDIN1(23) => ramainput_23_port, RAMDIN1(22) => 
                           ramainput_22_port, RAMDIN1(21) => ramainput_21_port,
                           RAMDIN1(20) => ramainput_20_port, RAMDIN1(19) => 
                           ramainput_19_port, RAMDIN1(18) => ramainput_18_port,
                           RAMDIN1(17) => ramainput_17_port, RAMDIN1(16) => 
                           ramainput_16_port, RAMDIN1(15) => ramainput_15_port,
                           RAMDIN1(14) => ramainput_14_port, RAMDIN1(13) => 
                           ramainput_13_port, RAMDIN1(12) => ramainput_12_port,
                           RAMDIN1(11) => ramainput_11_port, RAMDIN1(10) => 
                           ramainput_10_port, RAMDIN1(9) => ramainput_9_port, 
                           RAMDIN1(8) => ramainput_8_port, RAMDIN1(7) => 
                           ramainput_7_port, RAMDIN1(6) => ramainput_6_port, 
                           RAMDIN1(5) => ramainput_5_port, RAMDIN1(4) => 
                           ramainput_4_port, RAMDIN1(3) => ramainput_3_port, 
                           RAMDIN1(2) => ramainput_2_port, RAMDIN1(1) => 
                           ramainput_1_port, RAMDIN1(0) => ramainput_0_port, 
                           RAMDOUT1(127) => ramout1_127_port, RAMDOUT1(126) => 
                           ramout1_126_port, RAMDOUT1(125) => ramout1_125_port,
                           RAMDOUT1(124) => ramout1_124_port, RAMDOUT1(123) => 
                           ramout1_123_port, RAMDOUT1(122) => ramout1_122_port,
                           RAMDOUT1(121) => ramout1_121_port, RAMDOUT1(120) => 
                           ramout1_120_port, RAMDOUT1(119) => ramout1_119_port,
                           RAMDOUT1(118) => ramout1_118_port, RAMDOUT1(117) => 
                           ramout1_117_port, RAMDOUT1(116) => ramout1_116_port,
                           RAMDOUT1(115) => ramout1_115_port, RAMDOUT1(114) => 
                           ramout1_114_port, RAMDOUT1(113) => ramout1_113_port,
                           RAMDOUT1(112) => ramout1_112_port, RAMDOUT1(111) => 
                           ramout1_111_port, RAMDOUT1(110) => ramout1_110_port,
                           RAMDOUT1(109) => ramout1_109_port, RAMDOUT1(108) => 
                           ramout1_108_port, RAMDOUT1(107) => ramout1_107_port,
                           RAMDOUT1(106) => ramout1_106_port, RAMDOUT1(105) => 
                           ramout1_105_port, RAMDOUT1(104) => ramout1_104_port,
                           RAMDOUT1(103) => ramout1_103_port, RAMDOUT1(102) => 
                           ramout1_102_port, RAMDOUT1(101) => ramout1_101_port,
                           RAMDOUT1(100) => ramout1_100_port, RAMDOUT1(99) => 
                           ramout1_99_port, RAMDOUT1(98) => ramout1_98_port, 
                           RAMDOUT1(97) => ramout1_97_port, RAMDOUT1(96) => 
                           ramout1_96_port, RAMDOUT1(95) => ramout1_95_port, 
                           RAMDOUT1(94) => ramout1_94_port, RAMDOUT1(93) => 
                           ramout1_93_port, RAMDOUT1(92) => ramout1_92_port, 
                           RAMDOUT1(91) => ramout1_91_port, RAMDOUT1(90) => 
                           ramout1_90_port, RAMDOUT1(89) => ramout1_89_port, 
                           RAMDOUT1(88) => ramout1_88_port, RAMDOUT1(87) => 
                           ramout1_87_port, RAMDOUT1(86) => ramout1_86_port, 
                           RAMDOUT1(85) => ramout1_85_port, RAMDOUT1(84) => 
                           ramout1_84_port, RAMDOUT1(83) => ramout1_83_port, 
                           RAMDOUT1(82) => ramout1_82_port, RAMDOUT1(81) => 
                           ramout1_81_port, RAMDOUT1(80) => ramout1_80_port, 
                           RAMDOUT1(79) => ramout1_79_port, RAMDOUT1(78) => 
                           ramout1_78_port, RAMDOUT1(77) => ramout1_77_port, 
                           RAMDOUT1(76) => ramout1_76_port, RAMDOUT1(75) => 
                           ramout1_75_port, RAMDOUT1(74) => ramout1_74_port, 
                           RAMDOUT1(73) => ramout1_73_port, RAMDOUT1(72) => 
                           ramout1_72_port, RAMDOUT1(71) => ramout1_71_port, 
                           RAMDOUT1(70) => ramout1_70_port, RAMDOUT1(69) => 
                           ramout1_69_port, RAMDOUT1(68) => ramout1_68_port, 
                           RAMDOUT1(67) => ramout1_67_port, RAMDOUT1(66) => 
                           ramout1_66_port, RAMDOUT1(65) => ramout1_65_port, 
                           RAMDOUT1(64) => ramout1_64_port, RAMDOUT1(63) => 
                           ramout1_63_port, RAMDOUT1(62) => ramout1_62_port, 
                           RAMDOUT1(61) => ramout1_61_port, RAMDOUT1(60) => 
                           ramout1_60_port, RAMDOUT1(59) => ramout1_59_port, 
                           RAMDOUT1(58) => ramout1_58_port, RAMDOUT1(57) => 
                           ramout1_57_port, RAMDOUT1(56) => ramout1_56_port, 
                           RAMDOUT1(55) => ramout1_55_port, RAMDOUT1(54) => 
                           ramout1_54_port, RAMDOUT1(53) => ramout1_53_port, 
                           RAMDOUT1(52) => ramout1_52_port, RAMDOUT1(51) => 
                           ramout1_51_port, RAMDOUT1(50) => ramout1_50_port, 
                           RAMDOUT1(49) => ramout1_49_port, RAMDOUT1(48) => 
                           ramout1_48_port, RAMDOUT1(47) => ramout1_47_port, 
                           RAMDOUT1(46) => ramout1_46_port, RAMDOUT1(45) => 
                           ramout1_45_port, RAMDOUT1(44) => ramout1_44_port, 
                           RAMDOUT1(43) => ramout1_43_port, RAMDOUT1(42) => 
                           ramout1_42_port, RAMDOUT1(41) => ramout1_41_port, 
                           RAMDOUT1(40) => ramout1_40_port, RAMDOUT1(39) => 
                           ramout1_39_port, RAMDOUT1(38) => ramout1_38_port, 
                           RAMDOUT1(37) => ramout1_37_port, RAMDOUT1(36) => 
                           ramout1_36_port, RAMDOUT1(35) => ramout1_35_port, 
                           RAMDOUT1(34) => ramout1_34_port, RAMDOUT1(33) => 
                           ramout1_33_port, RAMDOUT1(32) => ramout1_32_port, 
                           RAMDOUT1(31) => ramout1_31_port, RAMDOUT1(30) => 
                           ramout1_30_port, RAMDOUT1(29) => ramout1_29_port, 
                           RAMDOUT1(28) => ramout1_28_port, RAMDOUT1(27) => 
                           ramout1_27_port, RAMDOUT1(26) => ramout1_26_port, 
                           RAMDOUT1(25) => ramout1_25_port, RAMDOUT1(24) => 
                           ramout1_24_port, RAMDOUT1(23) => ramout1_23_port, 
                           RAMDOUT1(22) => ramout1_22_port, RAMDOUT1(21) => 
                           ramout1_21_port, RAMDOUT1(20) => ramout1_20_port, 
                           RAMDOUT1(19) => ramout1_19_port, RAMDOUT1(18) => 
                           ramout1_18_port, RAMDOUT1(17) => ramout1_17_port, 
                           RAMDOUT1(16) => ramout1_16_port, RAMDOUT1(15) => 
                           ramout1_15_port, RAMDOUT1(14) => ramout1_14_port, 
                           RAMDOUT1(13) => ramout1_13_port, RAMDOUT1(12) => 
                           ramout1_12_port, RAMDOUT1(11) => ramout1_11_port, 
                           RAMDOUT1(10) => ramout1_10_port, RAMDOUT1(9) => 
                           ramout1_9_port, RAMDOUT1(8) => ramout1_8_port, 
                           RAMDOUT1(7) => ramout1_7_port, RAMDOUT1(6) => 
                           ramout1_6_port, RAMDOUT1(5) => ramout1_5_port, 
                           RAMDOUT1(4) => ramout1_4_port, RAMDOUT1(3) => 
                           ramout1_3_port, RAMDOUT1(2) => ramout1_2_port, 
                           RAMDOUT1(1) => ramout1_1_port, RAMDOUT1(0) => 
                           ramout1_0_port, RAMDOUT2(127) => ramout2_127_port, 
                           RAMDOUT2(126) => ramout2_126_port, RAMDOUT2(125) => 
                           ramout2_125_port, RAMDOUT2(124) => ramout2_124_port,
                           RAMDOUT2(123) => ramout2_123_port, RAMDOUT2(122) => 
                           ramout2_122_port, RAMDOUT2(121) => ramout2_121_port,
                           RAMDOUT2(120) => ramout2_120_port, RAMDOUT2(119) => 
                           ramout2_119_port, RAMDOUT2(118) => ramout2_118_port,
                           RAMDOUT2(117) => ramout2_117_port, RAMDOUT2(116) => 
                           ramout2_116_port, RAMDOUT2(115) => ramout2_115_port,
                           RAMDOUT2(114) => ramout2_114_port, RAMDOUT2(113) => 
                           ramout2_113_port, RAMDOUT2(112) => ramout2_112_port,
                           RAMDOUT2(111) => ramout2_111_port, RAMDOUT2(110) => 
                           ramout2_110_port, RAMDOUT2(109) => ramout2_109_port,
                           RAMDOUT2(108) => ramout2_108_port, RAMDOUT2(107) => 
                           ramout2_107_port, RAMDOUT2(106) => ramout2_106_port,
                           RAMDOUT2(105) => ramout2_105_port, RAMDOUT2(104) => 
                           ramout2_104_port, RAMDOUT2(103) => ramout2_103_port,
                           RAMDOUT2(102) => ramout2_102_port, RAMDOUT2(101) => 
                           ramout2_101_port, RAMDOUT2(100) => ramout2_100_port,
                           RAMDOUT2(99) => ramout2_99_port, RAMDOUT2(98) => 
                           ramout2_98_port, RAMDOUT2(97) => ramout2_97_port, 
                           RAMDOUT2(96) => ramout2_96_port, RAMDOUT2(95) => 
                           ramout2_95_port, RAMDOUT2(94) => ramout2_94_port, 
                           RAMDOUT2(93) => ramout2_93_port, RAMDOUT2(92) => 
                           ramout2_92_port, RAMDOUT2(91) => ramout2_91_port, 
                           RAMDOUT2(90) => ramout2_90_port, RAMDOUT2(89) => 
                           ramout2_89_port, RAMDOUT2(88) => ramout2_88_port, 
                           RAMDOUT2(87) => ramout2_87_port, RAMDOUT2(86) => 
                           ramout2_86_port, RAMDOUT2(85) => ramout2_85_port, 
                           RAMDOUT2(84) => ramout2_84_port, RAMDOUT2(83) => 
                           ramout2_83_port, RAMDOUT2(82) => ramout2_82_port, 
                           RAMDOUT2(81) => ramout2_81_port, RAMDOUT2(80) => 
                           ramout2_80_port, RAMDOUT2(79) => ramout2_79_port, 
                           RAMDOUT2(78) => ramout2_78_port, RAMDOUT2(77) => 
                           ramout2_77_port, RAMDOUT2(76) => ramout2_76_port, 
                           RAMDOUT2(75) => ramout2_75_port, RAMDOUT2(74) => 
                           ramout2_74_port, RAMDOUT2(73) => ramout2_73_port, 
                           RAMDOUT2(72) => ramout2_72_port, RAMDOUT2(71) => 
                           ramout2_71_port, RAMDOUT2(70) => ramout2_70_port, 
                           RAMDOUT2(69) => ramout2_69_port, RAMDOUT2(68) => 
                           ramout2_68_port, RAMDOUT2(67) => ramout2_67_port, 
                           RAMDOUT2(66) => ramout2_66_port, RAMDOUT2(65) => 
                           ramout2_65_port, RAMDOUT2(64) => ramout2_64_port, 
                           RAMDOUT2(63) => ramout2_63_port, RAMDOUT2(62) => 
                           ramout2_62_port, RAMDOUT2(61) => ramout2_61_port, 
                           RAMDOUT2(60) => ramout2_60_port, RAMDOUT2(59) => 
                           ramout2_59_port, RAMDOUT2(58) => ramout2_58_port, 
                           RAMDOUT2(57) => ramout2_57_port, RAMDOUT2(56) => 
                           ramout2_56_port, RAMDOUT2(55) => ramout2_55_port, 
                           RAMDOUT2(54) => ramout2_54_port, RAMDOUT2(53) => 
                           ramout2_53_port, RAMDOUT2(52) => ramout2_52_port, 
                           RAMDOUT2(51) => ramout2_51_port, RAMDOUT2(50) => 
                           ramout2_50_port, RAMDOUT2(49) => ramout2_49_port, 
                           RAMDOUT2(48) => ramout2_48_port, RAMDOUT2(47) => 
                           ramout2_47_port, RAMDOUT2(46) => ramout2_46_port, 
                           RAMDOUT2(45) => ramout2_45_port, RAMDOUT2(44) => 
                           ramout2_44_port, RAMDOUT2(43) => ramout2_43_port, 
                           RAMDOUT2(42) => ramout2_42_port, RAMDOUT2(41) => 
                           ramout2_41_port, RAMDOUT2(40) => ramout2_40_port, 
                           RAMDOUT2(39) => ramout2_39_port, RAMDOUT2(38) => 
                           ramout2_38_port, RAMDOUT2(37) => ramout2_37_port, 
                           RAMDOUT2(36) => ramout2_36_port, RAMDOUT2(35) => 
                           ramout2_35_port, RAMDOUT2(34) => ramout2_34_port, 
                           RAMDOUT2(33) => ramout2_33_port, RAMDOUT2(32) => 
                           ramout2_32_port, RAMDOUT2(31) => ramout2_31_port, 
                           RAMDOUT2(30) => ramout2_30_port, RAMDOUT2(29) => 
                           ramout2_29_port, RAMDOUT2(28) => ramout2_28_port, 
                           RAMDOUT2(27) => ramout2_27_port, RAMDOUT2(26) => 
                           ramout2_26_port, RAMDOUT2(25) => ramout2_25_port, 
                           RAMDOUT2(24) => ramout2_24_port, RAMDOUT2(23) => 
                           ramout2_23_port, RAMDOUT2(22) => ramout2_22_port, 
                           RAMDOUT2(21) => ramout2_21_port, RAMDOUT2(20) => 
                           ramout2_20_port, RAMDOUT2(19) => ramout2_19_port, 
                           RAMDOUT2(18) => ramout2_18_port, RAMDOUT2(17) => 
                           ramout2_17_port, RAMDOUT2(16) => ramout2_16_port, 
                           RAMDOUT2(15) => ramout2_15_port, RAMDOUT2(14) => 
                           ramout2_14_port, RAMDOUT2(13) => ramout2_13_port, 
                           RAMDOUT2(12) => ramout2_12_port, RAMDOUT2(11) => 
                           ramout2_11_port, RAMDOUT2(10) => ramout2_10_port, 
                           RAMDOUT2(9) => ramout2_9_port, RAMDOUT2(8) => 
                           ramout2_8_port, RAMDOUT2(7) => ramout2_7_port, 
                           RAMDOUT2(6) => ramout2_6_port, RAMDOUT2(5) => 
                           ramout2_5_port, RAMDOUT2(4) => ramout2_4_port, 
                           RAMDOUT2(3) => ramout2_3_port, RAMDOUT2(2) => 
                           ramout2_2_port, RAMDOUT2(1) => ramout2_1_port, 
                           RAMDOUT2(0) => ramout2_0_port, RAMWRITE1 => ramwrite
                           , clk => n40);
   XOODOO_PERM : 
                           xoodoo_round_ADDRESS_LEN128_ADDRESS_ENTRIES16_ADDRESS_ENTRIES_BITs4_1 
                           port map( RAMA(127) => ramout1_127_port, RAMA(126) 
                           => ramout1_126_port, RAMA(125) => ramout1_125_port, 
                           RAMA(124) => ramout1_124_port, RAMA(123) => 
                           ramout1_123_port, RAMA(122) => ramout1_122_port, 
                           RAMA(121) => ramout1_121_port, RAMA(120) => 
                           ramout1_120_port, RAMA(119) => ramout1_119_port, 
                           RAMA(118) => ramout1_118_port, RAMA(117) => 
                           ramout1_117_port, RAMA(116) => ramout1_116_port, 
                           RAMA(115) => ramout1_115_port, RAMA(114) => 
                           ramout1_114_port, RAMA(113) => ramout1_113_port, 
                           RAMA(112) => ramout1_112_port, RAMA(111) => 
                           ramout1_111_port, RAMA(110) => ramout1_110_port, 
                           RAMA(109) => ramout1_109_port, RAMA(108) => 
                           ramout1_108_port, RAMA(107) => ramout1_107_port, 
                           RAMA(106) => ramout1_106_port, RAMA(105) => 
                           ramout1_105_port, RAMA(104) => ramout1_104_port, 
                           RAMA(103) => ramout1_103_port, RAMA(102) => 
                           ramout1_102_port, RAMA(101) => ramout1_101_port, 
                           RAMA(100) => ramout1_100_port, RAMA(99) => 
                           ramout1_99_port, RAMA(98) => ramout1_98_port, 
                           RAMA(97) => ramout1_97_port, RAMA(96) => 
                           ramout1_96_port, RAMA(95) => ramout1_95_port, 
                           RAMA(94) => ramout1_94_port, RAMA(93) => 
                           ramout1_93_port, RAMA(92) => ramout1_92_port, 
                           RAMA(91) => ramout1_91_port, RAMA(90) => 
                           ramout1_90_port, RAMA(89) => ramout1_89_port, 
                           RAMA(88) => ramout1_88_port, RAMA(87) => 
                           ramout1_87_port, RAMA(86) => ramout1_86_port, 
                           RAMA(85) => ramout1_85_port, RAMA(84) => 
                           ramout1_84_port, RAMA(83) => ramout1_83_port, 
                           RAMA(82) => ramout1_82_port, RAMA(81) => 
                           ramout1_81_port, RAMA(80) => ramout1_80_port, 
                           RAMA(79) => ramout1_79_port, RAMA(78) => 
                           ramout1_78_port, RAMA(77) => ramout1_77_port, 
                           RAMA(76) => ramout1_76_port, RAMA(75) => 
                           ramout1_75_port, RAMA(74) => ramout1_74_port, 
                           RAMA(73) => ramout1_73_port, RAMA(72) => 
                           ramout1_72_port, RAMA(71) => ramout1_71_port, 
                           RAMA(70) => ramout1_70_port, RAMA(69) => 
                           ramout1_69_port, RAMA(68) => ramout1_68_port, 
                           RAMA(67) => ramout1_67_port, RAMA(66) => 
                           ramout1_66_port, RAMA(65) => ramout1_65_port, 
                           RAMA(64) => ramout1_64_port, RAMA(63) => 
                           ramout1_63_port, RAMA(62) => ramout1_62_port, 
                           RAMA(61) => ramout1_61_port, RAMA(60) => 
                           ramout1_60_port, RAMA(59) => ramout1_59_port, 
                           RAMA(58) => ramout1_58_port, RAMA(57) => 
                           ramout1_57_port, RAMA(56) => ramout1_56_port, 
                           RAMA(55) => ramout1_55_port, RAMA(54) => 
                           ramout1_54_port, RAMA(53) => ramout1_53_port, 
                           RAMA(52) => ramout1_52_port, RAMA(51) => 
                           ramout1_51_port, RAMA(50) => ramout1_50_port, 
                           RAMA(49) => ramout1_49_port, RAMA(48) => 
                           ramout1_48_port, RAMA(47) => ramout1_47_port, 
                           RAMA(46) => ramout1_46_port, RAMA(45) => 
                           ramout1_45_port, RAMA(44) => ramout1_44_port, 
                           RAMA(43) => ramout1_43_port, RAMA(42) => 
                           ramout1_42_port, RAMA(41) => ramout1_41_port, 
                           RAMA(40) => ramout1_40_port, RAMA(39) => 
                           ramout1_39_port, RAMA(38) => ramout1_38_port, 
                           RAMA(37) => ramout1_37_port, RAMA(36) => 
                           ramout1_36_port, RAMA(35) => ramout1_35_port, 
                           RAMA(34) => ramout1_34_port, RAMA(33) => 
                           ramout1_33_port, RAMA(32) => ramout1_32_port, 
                           RAMA(31) => ramout1_31_port, RAMA(30) => 
                           ramout1_30_port, RAMA(29) => ramout1_29_port, 
                           RAMA(28) => ramout1_28_port, RAMA(27) => 
                           ramout1_27_port, RAMA(26) => ramout1_26_port, 
                           RAMA(25) => ramout1_25_port, RAMA(24) => 
                           ramout1_24_port, RAMA(23) => ramout1_23_port, 
                           RAMA(22) => ramout1_22_port, RAMA(21) => 
                           ramout1_21_port, RAMA(20) => ramout1_20_port, 
                           RAMA(19) => ramout1_19_port, RAMA(18) => 
                           ramout1_18_port, RAMA(17) => ramout1_17_port, 
                           RAMA(16) => ramout1_16_port, RAMA(15) => 
                           ramout1_15_port, RAMA(14) => ramout1_14_port, 
                           RAMA(13) => ramout1_13_port, RAMA(12) => 
                           ramout1_12_port, RAMA(11) => ramout1_11_port, 
                           RAMA(10) => ramout1_10_port, RAMA(9) => 
                           ramout1_9_port, RAMA(8) => ramout1_8_port, RAMA(7) 
                           => ramout1_7_port, RAMA(6) => ramout1_6_port, 
                           RAMA(5) => ramout1_5_port, RAMA(4) => ramout1_4_port
                           , RAMA(3) => ramout1_3_port, RAMA(2) => 
                           ramout1_2_port, RAMA(1) => ramout1_1_port, RAMA(0) 
                           => ramout1_0_port, RAMB(127) => ramout2_127_port, 
                           RAMB(126) => ramout2_126_port, RAMB(125) => 
                           ramout2_125_port, RAMB(124) => ramout2_124_port, 
                           RAMB(123) => ramout2_123_port, RAMB(122) => 
                           ramout2_122_port, RAMB(121) => ramout2_121_port, 
                           RAMB(120) => ramout2_120_port, RAMB(119) => 
                           ramout2_119_port, RAMB(118) => ramout2_118_port, 
                           RAMB(117) => ramout2_117_port, RAMB(116) => 
                           ramout2_116_port, RAMB(115) => ramout2_115_port, 
                           RAMB(114) => ramout2_114_port, RAMB(113) => 
                           ramout2_113_port, RAMB(112) => ramout2_112_port, 
                           RAMB(111) => ramout2_111_port, RAMB(110) => 
                           ramout2_110_port, RAMB(109) => ramout2_109_port, 
                           RAMB(108) => ramout2_108_port, RAMB(107) => 
                           ramout2_107_port, RAMB(106) => ramout2_106_port, 
                           RAMB(105) => ramout2_105_port, RAMB(104) => 
                           ramout2_104_port, RAMB(103) => ramout2_103_port, 
                           RAMB(102) => ramout2_102_port, RAMB(101) => 
                           ramout2_101_port, RAMB(100) => ramout2_100_port, 
                           RAMB(99) => ramout2_99_port, RAMB(98) => 
                           ramout2_98_port, RAMB(97) => ramout2_97_port, 
                           RAMB(96) => ramout2_96_port, RAMB(95) => 
                           ramout2_95_port, RAMB(94) => ramout2_94_port, 
                           RAMB(93) => ramout2_93_port, RAMB(92) => 
                           ramout2_92_port, RAMB(91) => ramout2_91_port, 
                           RAMB(90) => ramout2_90_port, RAMB(89) => 
                           ramout2_89_port, RAMB(88) => ramout2_88_port, 
                           RAMB(87) => ramout2_87_port, RAMB(86) => 
                           ramout2_86_port, RAMB(85) => ramout2_85_port, 
                           RAMB(84) => ramout2_84_port, RAMB(83) => 
                           ramout2_83_port, RAMB(82) => ramout2_82_port, 
                           RAMB(81) => ramout2_81_port, RAMB(80) => 
                           ramout2_80_port, RAMB(79) => ramout2_79_port, 
                           RAMB(78) => ramout2_78_port, RAMB(77) => 
                           ramout2_77_port, RAMB(76) => ramout2_76_port, 
                           RAMB(75) => ramout2_75_port, RAMB(74) => 
                           ramout2_74_port, RAMB(73) => ramout2_73_port, 
                           RAMB(72) => ramout2_72_port, RAMB(71) => 
                           ramout2_71_port, RAMB(70) => ramout2_70_port, 
                           RAMB(69) => ramout2_69_port, RAMB(68) => 
                           ramout2_68_port, RAMB(67) => ramout2_67_port, 
                           RAMB(66) => ramout2_66_port, RAMB(65) => 
                           ramout2_65_port, RAMB(64) => ramout2_64_port, 
                           RAMB(63) => ramout2_63_port, RAMB(62) => 
                           ramout2_62_port, RAMB(61) => ramout2_61_port, 
                           RAMB(60) => ramout2_60_port, RAMB(59) => 
                           ramout2_59_port, RAMB(58) => ramout2_58_port, 
                           RAMB(57) => ramout2_57_port, RAMB(56) => 
                           ramout2_56_port, RAMB(55) => ramout2_55_port, 
                           RAMB(54) => ramout2_54_port, RAMB(53) => 
                           ramout2_53_port, RAMB(52) => ramout2_52_port, 
                           RAMB(51) => ramout2_51_port, RAMB(50) => 
                           ramout2_50_port, RAMB(49) => ramout2_49_port, 
                           RAMB(48) => ramout2_48_port, RAMB(47) => 
                           ramout2_47_port, RAMB(46) => ramout2_46_port, 
                           RAMB(45) => ramout2_45_port, RAMB(44) => 
                           ramout2_44_port, RAMB(43) => ramout2_43_port, 
                           RAMB(42) => ramout2_42_port, RAMB(41) => 
                           ramout2_41_port, RAMB(40) => ramout2_40_port, 
                           RAMB(39) => ramout2_39_port, RAMB(38) => 
                           ramout2_38_port, RAMB(37) => ramout2_37_port, 
                           RAMB(36) => ramout2_36_port, RAMB(35) => 
                           ramout2_35_port, RAMB(34) => ramout2_34_port, 
                           RAMB(33) => ramout2_33_port, RAMB(32) => 
                           ramout2_32_port, RAMB(31) => ramout2_31_port, 
                           RAMB(30) => ramout2_30_port, RAMB(29) => 
                           ramout2_29_port, RAMB(28) => ramout2_28_port, 
                           RAMB(27) => ramout2_27_port, RAMB(26) => 
                           ramout2_26_port, RAMB(25) => ramout2_25_port, 
                           RAMB(24) => ramout2_24_port, RAMB(23) => 
                           ramout2_23_port, RAMB(22) => ramout2_22_port, 
                           RAMB(21) => ramout2_21_port, RAMB(20) => 
                           ramout2_20_port, RAMB(19) => ramout2_19_port, 
                           RAMB(18) => ramout2_18_port, RAMB(17) => 
                           ramout2_17_port, RAMB(16) => ramout2_16_port, 
                           RAMB(15) => ramout2_15_port, RAMB(14) => 
                           ramout2_14_port, RAMB(13) => ramout2_13_port, 
                           RAMB(12) => ramout2_12_port, RAMB(11) => 
                           ramout2_11_port, RAMB(10) => ramout2_10_port, 
                           RAMB(9) => ramout2_9_port, RAMB(8) => ramout2_8_port
                           , RAMB(7) => ramout2_7_port, RAMB(6) => 
                           ramout2_6_port, RAMB(5) => ramout2_5_port, RAMB(4) 
                           => ramout2_4_port, RAMB(3) => ramout2_3_port, 
                           RAMB(2) => ramout2_2_port, RAMB(1) => ramout2_1_port
                           , RAMB(0) => ramout2_0_port, perm_output(127) => 
                           perm_output_127_port, perm_output(126) => 
                           perm_output_126_port, perm_output(125) => 
                           perm_output_125_port, perm_output(124) => 
                           perm_output_124_port, perm_output(123) => 
                           perm_output_123_port, perm_output(122) => 
                           perm_output_122_port, perm_output(121) => 
                           perm_output_121_port, perm_output(120) => 
                           perm_output_120_port, perm_output(119) => 
                           perm_output_119_port, perm_output(118) => 
                           perm_output_118_port, perm_output(117) => 
                           perm_output_117_port, perm_output(116) => 
                           perm_output_116_port, perm_output(115) => 
                           perm_output_115_port, perm_output(114) => 
                           perm_output_114_port, perm_output(113) => 
                           perm_output_113_port, perm_output(112) => 
                           perm_output_112_port, perm_output(111) => 
                           perm_output_111_port, perm_output(110) => 
                           perm_output_110_port, perm_output(109) => 
                           perm_output_109_port, perm_output(108) => 
                           perm_output_108_port, perm_output(107) => 
                           perm_output_107_port, perm_output(106) => 
                           perm_output_106_port, perm_output(105) => 
                           perm_output_105_port, perm_output(104) => 
                           perm_output_104_port, perm_output(103) => 
                           perm_output_103_port, perm_output(102) => 
                           perm_output_102_port, perm_output(101) => 
                           perm_output_101_port, perm_output(100) => 
                           perm_output_100_port, perm_output(99) => 
                           perm_output_99_port, perm_output(98) => 
                           perm_output_98_port, perm_output(97) => 
                           perm_output_97_port, perm_output(96) => 
                           perm_output_96_port, perm_output(95) => 
                           perm_output_95_port, perm_output(94) => 
                           perm_output_94_port, perm_output(93) => 
                           perm_output_93_port, perm_output(92) => 
                           perm_output_92_port, perm_output(91) => 
                           perm_output_91_port, perm_output(90) => 
                           perm_output_90_port, perm_output(89) => 
                           perm_output_89_port, perm_output(88) => 
                           perm_output_88_port, perm_output(87) => 
                           perm_output_87_port, perm_output(86) => 
                           perm_output_86_port, perm_output(85) => 
                           perm_output_85_port, perm_output(84) => 
                           perm_output_84_port, perm_output(83) => 
                           perm_output_83_port, perm_output(82) => 
                           perm_output_82_port, perm_output(81) => 
                           perm_output_81_port, perm_output(80) => 
                           perm_output_80_port, perm_output(79) => 
                           perm_output_79_port, perm_output(78) => 
                           perm_output_78_port, perm_output(77) => 
                           perm_output_77_port, perm_output(76) => 
                           perm_output_76_port, perm_output(75) => 
                           perm_output_75_port, perm_output(74) => 
                           perm_output_74_port, perm_output(73) => 
                           perm_output_73_port, perm_output(72) => 
                           perm_output_72_port, perm_output(71) => 
                           perm_output_71_port, perm_output(70) => 
                           perm_output_70_port, perm_output(69) => 
                           perm_output_69_port, perm_output(68) => 
                           perm_output_68_port, perm_output(67) => 
                           perm_output_67_port, perm_output(66) => 
                           perm_output_66_port, perm_output(65) => 
                           perm_output_65_port, perm_output(64) => 
                           perm_output_64_port, perm_output(63) => 
                           perm_output_63_port, perm_output(62) => 
                           perm_output_62_port, perm_output(61) => 
                           perm_output_61_port, perm_output(60) => 
                           perm_output_60_port, perm_output(59) => 
                           perm_output_59_port, perm_output(58) => 
                           perm_output_58_port, perm_output(57) => 
                           perm_output_57_port, perm_output(56) => 
                           perm_output_56_port, perm_output(55) => 
                           perm_output_55_port, perm_output(54) => 
                           perm_output_54_port, perm_output(53) => 
                           perm_output_53_port, perm_output(52) => 
                           perm_output_52_port, perm_output(51) => 
                           perm_output_51_port, perm_output(50) => 
                           perm_output_50_port, perm_output(49) => 
                           perm_output_49_port, perm_output(48) => 
                           perm_output_48_port, perm_output(47) => 
                           perm_output_47_port, perm_output(46) => 
                           perm_output_46_port, perm_output(45) => 
                           perm_output_45_port, perm_output(44) => 
                           perm_output_44_port, perm_output(43) => 
                           perm_output_43_port, perm_output(42) => 
                           perm_output_42_port, perm_output(41) => 
                           perm_output_41_port, perm_output(40) => 
                           perm_output_40_port, perm_output(39) => 
                           perm_output_39_port, perm_output(38) => 
                           perm_output_38_port, perm_output(37) => 
                           perm_output_37_port, perm_output(36) => 
                           perm_output_36_port, perm_output(35) => 
                           perm_output_35_port, perm_output(34) => 
                           perm_output_34_port, perm_output(33) => 
                           perm_output_33_port, perm_output(32) => 
                           perm_output_32_port, perm_output(31) => 
                           perm_output_31_port, perm_output(30) => 
                           perm_output_30_port, perm_output(29) => 
                           perm_output_29_port, perm_output(28) => 
                           perm_output_28_port, perm_output(27) => 
                           perm_output_27_port, perm_output(26) => 
                           perm_output_26_port, perm_output(25) => 
                           perm_output_25_port, perm_output(24) => 
                           perm_output_24_port, perm_output(23) => 
                           perm_output_23_port, perm_output(22) => 
                           perm_output_22_port, perm_output(21) => 
                           perm_output_21_port, perm_output(20) => 
                           perm_output_20_port, perm_output(19) => 
                           perm_output_19_port, perm_output(18) => 
                           perm_output_18_port, perm_output(17) => 
                           perm_output_17_port, perm_output(16) => 
                           perm_output_16_port, perm_output(15) => 
                           perm_output_15_port, perm_output(14) => 
                           perm_output_14_port, perm_output(13) => 
                           perm_output_13_port, perm_output(12) => 
                           perm_output_12_port, perm_output(11) => 
                           perm_output_11_port, perm_output(10) => 
                           perm_output_10_port, perm_output(9) => 
                           perm_output_9_port, perm_output(8) => 
                           perm_output_8_port, perm_output(7) => 
                           perm_output_7_port, perm_output(6) => 
                           perm_output_6_port, perm_output(5) => 
                           perm_output_5_port, perm_output(4) => 
                           perm_output_4_port, perm_output(3) => 
                           perm_output_3_port, perm_output(2) => 
                           perm_output_2_port, perm_output(1) => 
                           perm_output_1_port, perm_output(0) => 
                           perm_output_0_port, ADDRA(3) => perm_addr_3_port, 
                           ADDRA(2) => perm_addr_2_port, ADDRA(1) => 
                           perm_addr_1_port, ADDRA(0) => perm_addr_0_port, 
                           ADDRB(3) => perm_addr2_3_port, ADDRB(2) => 
                           perm_addr2_2_port, ADDRB(1) => perm_addr2_1_port, 
                           ADDRB(0) => perm_addr2_0_port, RNDCTR(3) => 
                           rnd_counter_3_port, RNDCTR(2) => rnd_counter_2_port,
                           RNDCTR(1) => rnd_counter_1_port, RNDCTR(0) => 
                           rnd_counter_0_port, ins_counter(4) => 
                           ins_counter_4_port, ins_counter(3) => 
                           ins_counter_3_port, ins_counter(2) => 
                           ins_counter_2_port, ins_counter(1) => 
                           ins_counter_1_port, ins_counter(0) => 
                           ins_counter_0_port);
   round_counter : counter_num_bits4_1_0 port map( clk => n40, load => load_rnd
                           , enable => en_rnd, start_value(3) => X_Logic0_port,
                           start_value(2) => X_Logic0_port, start_value(1) => 
                           X_Logic0_port, start_value(0) => X_Logic0_port, q(3)
                           => rnd_counter_3_port, q(2) => rnd_counter_2_port, 
                           q(1) => rnd_counter_1_port, q(0) => 
                           rnd_counter_0_port);
   E_ins_counter : counter_num_bits5_1 port map( clk => n40, load => load_ins, 
                           enable => n62, start_value(4) => 
                           ins_start_value_4_port, start_value(3) => 
                           ins_start_value_3_port, start_value(2) => 
                           ins_start_value_0, start_value(1) => X_Logic0_port, 
                           start_value(0) => ins_start_value_0, q(4) => 
                           ins_counter_4_port, q(3) => ins_counter_3_port, q(2)
                           => ins_counter_2_port, q(1) => ins_counter_1_port, 
                           q(0) => ins_counter_0_port);
   E_dcount : counter_num_bits4_1_1 port map( clk => n40, load => load_dcount, 
                           enable => en_dcount, start_value(3) => 
                           dcount_start_value_3, start_value(2) => 
                           X_Logic0_port, start_value(1) => 
                           dcount_start_value_3, start_value(0) => 
                           dcount_start_value_3, q(3) => dcount_3_port, q(2) =>
                           dcount_2_port, q(1) => dcount_1_port, q(0) => 
                           dcount_0_port);
   cyc_ops : cyclist_ops_RAM_LEN128_DATA_LEN32_1 port map( 
                           cyc_state_update_sel(1) => 
                           cyc_state_update_sel_1_port, cyc_state_update_sel(0)
                           => cyc_state_update_sel_0_port, xor_sel(1) => 
                           xor_sel_1_port, xor_sel(0) => n247, cycd_sel(1) => 
                           cycd_sel_1_port, cycd_sel(0) => cycd_sel_0_port, 
                           extract_sel => extract_sel, addr_sel2 => 
                           addr_sel_1_port, ramoutd1(127) => ramout1_127_port, 
                           ramoutd1(126) => ramout1_126_port, ramoutd1(125) => 
                           ramout1_125_port, ramoutd1(124) => ramout1_124_port,
                           ramoutd1(123) => ramout1_123_port, ramoutd1(122) => 
                           ramout1_122_port, ramoutd1(121) => ramout1_121_port,
                           ramoutd1(120) => ramout1_120_port, ramoutd1(119) => 
                           ramout1_119_port, ramoutd1(118) => ramout1_118_port,
                           ramoutd1(117) => ramout1_117_port, ramoutd1(116) => 
                           ramout1_116_port, ramoutd1(115) => ramout1_115_port,
                           ramoutd1(114) => ramout1_114_port, ramoutd1(113) => 
                           ramout1_113_port, ramoutd1(112) => ramout1_112_port,
                           ramoutd1(111) => ramout1_111_port, ramoutd1(110) => 
                           ramout1_110_port, ramoutd1(109) => ramout1_109_port,
                           ramoutd1(108) => ramout1_108_port, ramoutd1(107) => 
                           ramout1_107_port, ramoutd1(106) => ramout1_106_port,
                           ramoutd1(105) => ramout1_105_port, ramoutd1(104) => 
                           ramout1_104_port, ramoutd1(103) => ramout1_103_port,
                           ramoutd1(102) => ramout1_102_port, ramoutd1(101) => 
                           ramout1_101_port, ramoutd1(100) => ramout1_100_port,
                           ramoutd1(99) => ramout1_99_port, ramoutd1(98) => 
                           ramout1_98_port, ramoutd1(97) => ramout1_97_port, 
                           ramoutd1(96) => ramout1_96_port, ramoutd1(95) => 
                           ramout1_95_port, ramoutd1(94) => ramout1_94_port, 
                           ramoutd1(93) => ramout1_93_port, ramoutd1(92) => 
                           ramout1_92_port, ramoutd1(91) => ramout1_91_port, 
                           ramoutd1(90) => ramout1_90_port, ramoutd1(89) => 
                           ramout1_89_port, ramoutd1(88) => ramout1_88_port, 
                           ramoutd1(87) => ramout1_87_port, ramoutd1(86) => 
                           ramout1_86_port, ramoutd1(85) => ramout1_85_port, 
                           ramoutd1(84) => ramout1_84_port, ramoutd1(83) => 
                           ramout1_83_port, ramoutd1(82) => ramout1_82_port, 
                           ramoutd1(81) => ramout1_81_port, ramoutd1(80) => 
                           ramout1_80_port, ramoutd1(79) => ramout1_79_port, 
                           ramoutd1(78) => ramout1_78_port, ramoutd1(77) => 
                           ramout1_77_port, ramoutd1(76) => ramout1_76_port, 
                           ramoutd1(75) => ramout1_75_port, ramoutd1(74) => 
                           ramout1_74_port, ramoutd1(73) => ramout1_73_port, 
                           ramoutd1(72) => ramout1_72_port, ramoutd1(71) => 
                           ramout1_71_port, ramoutd1(70) => ramout1_70_port, 
                           ramoutd1(69) => ramout1_69_port, ramoutd1(68) => 
                           ramout1_68_port, ramoutd1(67) => ramout1_67_port, 
                           ramoutd1(66) => ramout1_66_port, ramoutd1(65) => 
                           ramout1_65_port, ramoutd1(64) => ramout1_64_port, 
                           ramoutd1(63) => ramout1_63_port, ramoutd1(62) => 
                           ramout1_62_port, ramoutd1(61) => ramout1_61_port, 
                           ramoutd1(60) => ramout1_60_port, ramoutd1(59) => 
                           ramout1_59_port, ramoutd1(58) => ramout1_58_port, 
                           ramoutd1(57) => ramout1_57_port, ramoutd1(56) => 
                           ramout1_56_port, ramoutd1(55) => ramout1_55_port, 
                           ramoutd1(54) => ramout1_54_port, ramoutd1(53) => 
                           ramout1_53_port, ramoutd1(52) => ramout1_52_port, 
                           ramoutd1(51) => ramout1_51_port, ramoutd1(50) => 
                           ramout1_50_port, ramoutd1(49) => ramout1_49_port, 
                           ramoutd1(48) => ramout1_48_port, ramoutd1(47) => 
                           ramout1_47_port, ramoutd1(46) => ramout1_46_port, 
                           ramoutd1(45) => ramout1_45_port, ramoutd1(44) => 
                           ramout1_44_port, ramoutd1(43) => ramout1_43_port, 
                           ramoutd1(42) => ramout1_42_port, ramoutd1(41) => 
                           ramout1_41_port, ramoutd1(40) => ramout1_40_port, 
                           ramoutd1(39) => ramout1_39_port, ramoutd1(38) => 
                           ramout1_38_port, ramoutd1(37) => ramout1_37_port, 
                           ramoutd1(36) => ramout1_36_port, ramoutd1(35) => 
                           ramout1_35_port, ramoutd1(34) => ramout1_34_port, 
                           ramoutd1(33) => ramout1_33_port, ramoutd1(32) => 
                           ramout1_32_port, ramoutd1(31) => ramout1_31_port, 
                           ramoutd1(30) => ramout1_30_port, ramoutd1(29) => 
                           ramout1_29_port, ramoutd1(28) => ramout1_28_port, 
                           ramoutd1(27) => ramout1_27_port, ramoutd1(26) => 
                           ramout1_26_port, ramoutd1(25) => ramout1_25_port, 
                           ramoutd1(24) => ramout1_24_port, ramoutd1(23) => 
                           ramout1_23_port, ramoutd1(22) => ramout1_22_port, 
                           ramoutd1(21) => ramout1_21_port, ramoutd1(20) => 
                           ramout1_20_port, ramoutd1(19) => ramout1_19_port, 
                           ramoutd1(18) => ramout1_18_port, ramoutd1(17) => 
                           ramout1_17_port, ramoutd1(16) => ramout1_16_port, 
                           ramoutd1(15) => ramout1_15_port, ramoutd1(14) => 
                           ramout1_14_port, ramoutd1(13) => ramout1_13_port, 
                           ramoutd1(12) => ramout1_12_port, ramoutd1(11) => 
                           ramout1_11_port, ramoutd1(10) => ramout1_10_port, 
                           ramoutd1(9) => ramout1_9_port, ramoutd1(8) => 
                           ramout1_8_port, ramoutd1(7) => ramout1_7_port, 
                           ramoutd1(6) => ramout1_6_port, ramoutd1(5) => 
                           ramout1_5_port, ramoutd1(4) => ramout1_4_port, 
                           ramoutd1(3) => ramout1_3_port, ramoutd1(2) => 
                           ramout1_2_port, ramoutd1(1) => ramout1_1_port, 
                           ramoutd1(0) => ramout1_0_port, key(31) => key(7), 
                           key(30) => key(6), key(29) => key(5), key(28) => 
                           key(4), key(27) => key(3), key(26) => key(2), 
                           key(25) => key(1), key(24) => key(0), key(23) => 
                           key(15), key(22) => key(14), key(21) => key(13), 
                           key(20) => key(12), key(19) => key(11), key(18) => 
                           key(10), key(17) => key(9), key(16) => key(8), 
                           key(15) => key(23), key(14) => key(22), key(13) => 
                           key(21), key(12) => key(20), key(11) => key(19), 
                           key(10) => key(18), key(9) => key(17), key(8) => 
                           key(16), key(7) => key(31), key(6) => key(30), 
                           key(5) => key(29), key(4) => key(28), key(3) => 
                           key(27), key(2) => key(26), key(1) => key(25), 
                           key(0) => key(24), bdi_data(31) => bdi(7), 
                           bdi_data(30) => bdi(6), bdi_data(29) => bdi(5), 
                           bdi_data(28) => bdi(4), bdi_data(27) => bdi(3), 
                           bdi_data(26) => bdi(2), bdi_data(25) => bdi(1), 
                           bdi_data(24) => bdi(0), bdi_data(23) => bdi(15), 
                           bdi_data(22) => bdi(14), bdi_data(21) => bdi(13), 
                           bdi_data(20) => bdi(12), bdi_data(19) => bdi(11), 
                           bdi_data(18) => bdi(10), bdi_data(17) => bdi(9), 
                           bdi_data(16) => bdi(8), bdi_data(15) => bdi(23), 
                           bdi_data(14) => bdi(22), bdi_data(13) => bdi(21), 
                           bdi_data(12) => bdi(20), bdi_data(11) => bdi(19), 
                           bdi_data(10) => bdi(18), bdi_data(9) => bdi(17), 
                           bdi_data(8) => bdi(16), bdi_data(7) => bdi(31), 
                           bdi_data(6) => bdi(30), bdi_data(5) => bdi(29), 
                           bdi_data(4) => bdi(28), bdi_data(3) => bdi(27), 
                           bdi_data(2) => bdi(26), bdi_data(1) => bdi(25), 
                           bdi_data(0) => bdi(24), cu_cd(7) => n255, cu_cd(6) 
                           => cu_cd_s_6_port, cu_cd(5) => X_Logic0_port, 
                           cu_cd(4) => X_Logic0_port, cu_cd(3) => X_Logic0_port
                           , cu_cd(2) => X_Logic0_port, cu_cd(1) => cu_cd_s_1, 
                           cu_cd(0) => n253, dcount_in(1) => dcount_1_port, 
                           dcount_in(0) => dcount_0_port, cyc_state_update(127)
                           => cyc_state_update_127_port, cyc_state_update(126) 
                           => cyc_state_update_126_port, cyc_state_update(125) 
                           => cyc_state_update_125_port, cyc_state_update(124) 
                           => cyc_state_update_124_port, cyc_state_update(123) 
                           => cyc_state_update_123_port, cyc_state_update(122) 
                           => cyc_state_update_122_port, cyc_state_update(121) 
                           => cyc_state_update_121_port, cyc_state_update(120) 
                           => cyc_state_update_120_port, cyc_state_update(119) 
                           => cyc_state_update_119_port, cyc_state_update(118) 
                           => cyc_state_update_118_port, cyc_state_update(117) 
                           => cyc_state_update_117_port, cyc_state_update(116) 
                           => cyc_state_update_116_port, cyc_state_update(115) 
                           => cyc_state_update_115_port, cyc_state_update(114) 
                           => cyc_state_update_114_port, cyc_state_update(113) 
                           => cyc_state_update_113_port, cyc_state_update(112) 
                           => cyc_state_update_112_port, cyc_state_update(111) 
                           => cyc_state_update_111_port, cyc_state_update(110) 
                           => cyc_state_update_110_port, cyc_state_update(109) 
                           => cyc_state_update_109_port, cyc_state_update(108) 
                           => cyc_state_update_108_port, cyc_state_update(107) 
                           => cyc_state_update_107_port, cyc_state_update(106) 
                           => cyc_state_update_106_port, cyc_state_update(105) 
                           => cyc_state_update_105_port, cyc_state_update(104) 
                           => cyc_state_update_104_port, cyc_state_update(103) 
                           => cyc_state_update_103_port, cyc_state_update(102) 
                           => cyc_state_update_102_port, cyc_state_update(101) 
                           => cyc_state_update_101_port, cyc_state_update(100) 
                           => cyc_state_update_100_port, cyc_state_update(99) 
                           => cyc_state_update_99_port, cyc_state_update(98) =>
                           cyc_state_update_98_port, cyc_state_update(97) => 
                           cyc_state_update_97_port, cyc_state_update(96) => 
                           cyc_state_update_96_port, cyc_state_update(95) => 
                           cyc_state_update_95_port, cyc_state_update(94) => 
                           cyc_state_update_94_port, cyc_state_update(93) => 
                           cyc_state_update_93_port, cyc_state_update(92) => 
                           cyc_state_update_92_port, cyc_state_update(91) => 
                           cyc_state_update_91_port, cyc_state_update(90) => 
                           cyc_state_update_90_port, cyc_state_update(89) => 
                           cyc_state_update_89_port, cyc_state_update(88) => 
                           cyc_state_update_88_port, cyc_state_update(87) => 
                           cyc_state_update_87_port, cyc_state_update(86) => 
                           cyc_state_update_86_port, cyc_state_update(85) => 
                           cyc_state_update_85_port, cyc_state_update(84) => 
                           cyc_state_update_84_port, cyc_state_update(83) => 
                           cyc_state_update_83_port, cyc_state_update(82) => 
                           cyc_state_update_82_port, cyc_state_update(81) => 
                           cyc_state_update_81_port, cyc_state_update(80) => 
                           cyc_state_update_80_port, cyc_state_update(79) => 
                           cyc_state_update_79_port, cyc_state_update(78) => 
                           cyc_state_update_78_port, cyc_state_update(77) => 
                           cyc_state_update_77_port, cyc_state_update(76) => 
                           cyc_state_update_76_port, cyc_state_update(75) => 
                           cyc_state_update_75_port, cyc_state_update(74) => 
                           cyc_state_update_74_port, cyc_state_update(73) => 
                           cyc_state_update_73_port, cyc_state_update(72) => 
                           cyc_state_update_72_port, cyc_state_update(71) => 
                           cyc_state_update_71_port, cyc_state_update(70) => 
                           cyc_state_update_70_port, cyc_state_update(69) => 
                           cyc_state_update_69_port, cyc_state_update(68) => 
                           cyc_state_update_68_port, cyc_state_update(67) => 
                           cyc_state_update_67_port, cyc_state_update(66) => 
                           cyc_state_update_66_port, cyc_state_update(65) => 
                           cyc_state_update_65_port, cyc_state_update(64) => 
                           cyc_state_update_64_port, cyc_state_update(63) => 
                           cyc_state_update_63_port, cyc_state_update(62) => 
                           cyc_state_update_62_port, cyc_state_update(61) => 
                           cyc_state_update_61_port, cyc_state_update(60) => 
                           cyc_state_update_60_port, cyc_state_update(59) => 
                           cyc_state_update_59_port, cyc_state_update(58) => 
                           cyc_state_update_58_port, cyc_state_update(57) => 
                           cyc_state_update_57_port, cyc_state_update(56) => 
                           cyc_state_update_56_port, cyc_state_update(55) => 
                           cyc_state_update_55_port, cyc_state_update(54) => 
                           cyc_state_update_54_port, cyc_state_update(53) => 
                           cyc_state_update_53_port, cyc_state_update(52) => 
                           cyc_state_update_52_port, cyc_state_update(51) => 
                           cyc_state_update_51_port, cyc_state_update(50) => 
                           cyc_state_update_50_port, cyc_state_update(49) => 
                           cyc_state_update_49_port, cyc_state_update(48) => 
                           cyc_state_update_48_port, cyc_state_update(47) => 
                           cyc_state_update_47_port, cyc_state_update(46) => 
                           cyc_state_update_46_port, cyc_state_update(45) => 
                           cyc_state_update_45_port, cyc_state_update(44) => 
                           cyc_state_update_44_port, cyc_state_update(43) => 
                           cyc_state_update_43_port, cyc_state_update(42) => 
                           cyc_state_update_42_port, cyc_state_update(41) => 
                           cyc_state_update_41_port, cyc_state_update(40) => 
                           cyc_state_update_40_port, cyc_state_update(39) => 
                           cyc_state_update_39_port, cyc_state_update(38) => 
                           cyc_state_update_38_port, cyc_state_update(37) => 
                           cyc_state_update_37_port, cyc_state_update(36) => 
                           cyc_state_update_36_port, cyc_state_update(35) => 
                           cyc_state_update_35_port, cyc_state_update(34) => 
                           cyc_state_update_34_port, cyc_state_update(33) => 
                           cyc_state_update_33_port, cyc_state_update(32) => 
                           cyc_state_update_32_port, cyc_state_update(31) => 
                           cyc_state_update_31_port, cyc_state_update(30) => 
                           cyc_state_update_30_port, cyc_state_update(29) => 
                           cyc_state_update_29_port, cyc_state_update(28) => 
                           cyc_state_update_28_port, cyc_state_update(27) => 
                           cyc_state_update_27_port, cyc_state_update(26) => 
                           cyc_state_update_26_port, cyc_state_update(25) => 
                           cyc_state_update_25_port, cyc_state_update(24) => 
                           cyc_state_update_24_port, cyc_state_update(23) => 
                           cyc_state_update_23_port, cyc_state_update(22) => 
                           cyc_state_update_22_port, cyc_state_update(21) => 
                           cyc_state_update_21_port, cyc_state_update(20) => 
                           cyc_state_update_20_port, cyc_state_update(19) => 
                           cyc_state_update_19_port, cyc_state_update(18) => 
                           cyc_state_update_18_port, cyc_state_update(17) => 
                           cyc_state_update_17_port, cyc_state_update(16) => 
                           cyc_state_update_16_port, cyc_state_update(15) => 
                           cyc_state_update_15_port, cyc_state_update(14) => 
                           cyc_state_update_14_port, cyc_state_update(13) => 
                           cyc_state_update_13_port, cyc_state_update(12) => 
                           cyc_state_update_12_port, cyc_state_update(11) => 
                           cyc_state_update_11_port, cyc_state_update(10) => 
                           cyc_state_update_10_port, cyc_state_update(9) => 
                           cyc_state_update_9_port, cyc_state_update(8) => 
                           cyc_state_update_8_port, cyc_state_update(7) => 
                           cyc_state_update_7_port, cyc_state_update(6) => 
                           cyc_state_update_6_port, cyc_state_update(5) => 
                           cyc_state_update_5_port, cyc_state_update(4) => 
                           cyc_state_update_4_port, cyc_state_update(3) => 
                           cyc_state_update_3_port, cyc_state_update(2) => 
                           cyc_state_update_2_port, cyc_state_update(1) => 
                           cyc_state_update_1_port, cyc_state_update(0) => 
                           cyc_state_update_0_port, bdo_out(31) => n267, 
                           bdo_out(30) => n268, bdo_out(29) => n269, 
                           bdo_out(28) => bdo_4_port, bdo_out(27) => n270, 
                           bdo_out(26) => bdo_2_port, bdo_out(25) => n271, 
                           bdo_out(24) => bdo_0_port, bdo_out(23) => 
                           bdo_15_port, bdo_out(22) => bdo_14_port, bdo_out(21)
                           => bdo_13_port, bdo_out(20) => bdo_12_port, 
                           bdo_out(19) => bdo_11_port, bdo_out(18) => 
                           bdo_10_port, bdo_out(17) => bdo_9_port, bdo_out(16) 
                           => bdo_8_port, bdo_out(15) => bdo_23_port, 
                           bdo_out(14) => bdo_22_port, bdo_out(13) => 
                           bdo_21_port, bdo_out(12) => bdo_20_port, bdo_out(11)
                           => bdo_19_port, bdo_out(10) => bdo_18_port, 
                           bdo_out(9) => bdo_17_port, bdo_out(8) => bdo_16_port
                           , bdo_out(7) => n265, bdo_out(6) => n266, bdo_out(5)
                           => bdo_29_port, bdo_out(4) => bdo_28_port, 
                           bdo_out(3) => bdo_27_port, bdo_out(2) => bdo_26_port
                           , bdo_out(1) => bdo_25_port, bdo_out(0) => 
                           bdo_24_port);
   r195 : CryptoCore_1_DW01_cmp6_0 port map( A(31) => bdi(7), A(30) => bdi(6), 
                           A(29) => bdi(5), A(28) => bdi(4), A(27) => bdi(3), 
                           A(26) => bdi(2), A(25) => bdi(1), A(24) => bdi(0), 
                           A(23) => bdi(15), A(22) => bdi(14), A(21) => bdi(13)
                           , A(20) => bdi(12), A(19) => bdi(11), A(18) => 
                           bdi(10), A(17) => bdi(9), A(16) => bdi(8), A(15) => 
                           bdi(23), A(14) => bdi(22), A(13) => bdi(21), A(12) 
                           => bdi(20), A(11) => bdi(19), A(10) => bdi(18), A(9)
                           => bdi(17), A(8) => bdi(16), A(7) => bdi(31), A(6) 
                           => bdi(30), A(5) => bdi(29), A(4) => bdi(28), A(3) 
                           => bdi(27), A(2) => bdi(26), A(1) => bdi(25), A(0) 
                           => bdi(24), B(31) => n267, B(30) => n268, B(29) => 
                           n269, B(28) => bdo_4_port, B(27) => n270, B(26) => 
                           bdo_2_port, B(25) => n271, B(24) => bdo_0_port, 
                           B(23) => bdo_15_port, B(22) => bdo_14_port, B(21) =>
                           bdo_13_port, B(20) => bdo_12_port, B(19) => 
                           bdo_11_port, B(18) => bdo_10_port, B(17) => 
                           bdo_9_port, B(16) => bdo_8_port, B(15) => 
                           bdo_23_port, B(14) => bdo_22_port, B(13) => 
                           bdo_21_port, B(12) => bdo_20_port, B(11) => 
                           bdo_19_port, B(10) => bdo_18_port, B(9) => 
                           bdo_17_port, B(8) => bdo_16_port, B(7) => n265, B(6)
                           => n266, B(5) => bdo_29_port, B(4) => bdo_28_port, 
                           B(3) => bdo_27_port, B(2) => bdo_26_port, B(1) => 
                           bdo_25_port, B(0) => bdo_24_port, TC => n1, LT => 
                           n_3226, GT => n_3227, EQ => n_3228, LE => n_3229, GE
                           => n_3230, NE => N275);
   cyc_s_reg_2_inst : DFFX1 port map( D => n212, CLK => n40, Q => cyc_s_2_port,
                           QN => n44);
   cyc_s_reg_1_inst : DFFX1 port map( D => n209, CLK => n40, Q => cyc_s_1_port,
                           QN => n45);
   U3 : AND2X4 port map( IN1 => n15, IN2 => perm_addr_3_port, Q => 
                           addrmux2_3_port);
   U5 : AND2X4 port map( IN1 => n147, IN2 => cyc_s_0_port, Q => n2);
   U6 : OR2X2 port map( IN1 => n35, IN2 => n32, Q => n159);
   U7 : AO22X2 port map( IN1 => perm_output_99_port, IN2 => n222, IN3 => 
                           cyc_state_update_99_port, IN4 => n47, Q => 
                           ramainput_99_port);
   U8 : AO22X1 port map( IN1 => perm_output_24_port, IN2 => n203, IN3 => 
                           cyc_state_update_24_port, IN4 => n57, Q => 
                           ramainput_24_port);
   U9 : AO22X1 port map( IN1 => perm_output_41_port, IN2 => n216, IN3 => 
                           cyc_state_update_41_port, IN4 => n56, Q => 
                           ramainput_41_port);
   U10 : AO22X2 port map( IN1 => perm_output_103_port, IN2 => n197, IN3 => 
                           cyc_state_update_103_port, IN4 => n61, Q => 
                           ramainput_103_port);
   U11 : AO221X2 port map( IN1 => perm_addr_1_port, IN2 => n16, IN3 => 
                           dcount_3_port, IN4 => n4, IN5 => addr_sel_1_port, Q 
                           => addrmux2_1_port);
   U12 : DELLN2X2 port map( INP => n11, Z => n37);
   U13 : DELLN1X2 port map( INP => n159, Z => n3);
   U14 : OR2X4 port map( IN1 => addr_sel_1_port, IN2 => n36, Q => 
                           xor_sel_1_port);
   U15 : AOI21X1 port map( IN1 => n2, IN2 => n7, IN3 => n36, QN => n64);
   U16 : IBUFFX16 port map( INP => n41, ZN => n251);
   U17 : NAND3X1 port map( IN1 => n81, IN2 => n159, IN3 => n156, QN => 
                           addr_sel_1_port);
   U18 : AND2X1 port map( IN1 => n15, IN2 => perm_addr_2_port, Q => 
                           addrmux2_2_port);
   U19 : AO221X1 port map( IN1 => n165, IN2 => n181, IN3 => n182, IN4 => n8, 
                           IN5 => bdo_type_3_port, Q => bdo_valid);
   U20 : AO22X1 port map( IN1 => n245, IN2 => calling_state_2_port, IN3 => n85,
                           IN4 => n251, Q => n207);
   U21 : NAND3X0 port map( IN1 => n248, IN2 => n251, IN3 => n132, QN => n131);
   U22 : NAND4X1 port map( IN1 => n157, IN2 => n81, IN3 => n64, IN4 => n6, QN 
                           => n4);
   U23 : AND2X1 port map( IN1 => n243, IN2 => n140, Q => n5);
   U24 : AO22X2 port map( IN1 => perm_output_43_port, IN2 => n216, IN3 => 
                           cyc_state_update_43_port, IN4 => n56, Q => 
                           ramainput_43_port);
   U25 : AO22X2 port map( IN1 => perm_output_22_port, IN2 => n203, IN3 => 
                           cyc_state_update_22_port, IN4 => n58, Q => 
                           ramainput_22_port);
   U26 : AO22X2 port map( IN1 => perm_output_48_port, IN2 => n203, IN3 => 
                           cyc_state_update_48_port, IN4 => n55, Q => 
                           ramainput_48_port);
   U27 : AO22X2 port map( IN1 => perm_output_5_port, IN2 => n218, IN3 => 
                           cyc_state_update_5_port, IN4 => n50, Q => 
                           ramainput_5_port);
   U28 : AO22X2 port map( IN1 => perm_output_101_port, IN2 => n197, IN3 => 
                           cyc_state_update_101_port, IN4 => n61, Q => 
                           ramainput_101_port);
   U29 : AO22X2 port map( IN1 => perm_output_107_port, IN2 => n200, IN3 => 
                           cyc_state_update_107_port, IN4 => n60, Q => 
                           ramainput_107_port);
   U30 : AO22X2 port map( IN1 => perm_output_3_port, IN2 => n215, IN3 => 
                           cyc_state_update_3_port, IN4 => n56, Q => 
                           ramainput_3_port);
   U31 : AO22X2 port map( IN1 => perm_output_113_port, IN2 => n201, IN3 => 
                           cyc_state_update_113_port, IN4 => n60, Q => 
                           ramainput_113_port);
   U32 : AO22X2 port map( IN1 => perm_output_76_port, IN2 => n220, IN3 => 
                           cyc_state_update_76_port, IN4 => n49, Q => 
                           ramainput_76_port);
   U33 : AND2X4 port map( IN1 => n101, IN2 => n68, Q => n6);
   U34 : AND2X1 port map( IN1 => n101, IN2 => n68, Q => n199);
   U35 : AO22X2 port map( IN1 => perm_output_124_port, IN2 => n200, IN3 => 
                           cyc_state_update_124_port, IN4 => n59, Q => 
                           ramainput_124_port);
   U36 : IBUFFX16 port map( INP => n36, ZN => n173);
   U37 : IBUFFX16 port map( INP => n162, ZN => n7);
   U38 : INVX0 port map( INP => N275, ZN => n229);
   U39 : DELLN2X2 port map( INP => n36, Z => n8);
   U40 : DELLN2X2 port map( INP => n101, Z => n9);
   U41 : AO22X2 port map( IN1 => perm_output_102_port, IN2 => n197, IN3 => 
                           cyc_state_update_102_port, IN4 => n61, Q => 
                           ramainput_102_port);
   U42 : NOR2X0 port map( IN1 => n35, IN2 => n162, QN => n10);
   U43 : NOR2X0 port map( IN1 => n10, IN2 => n36, QN => n11);
   U44 : AND4X1 port map( IN1 => n199, IN2 => n64, IN3 => n81, IN4 => n157, Q 
                           => n12);
   U45 : AND2X1 port map( IN1 => cyc_s_1_port, IN2 => cyc_s_2_port, Q => n148);
   U46 : NAND3X4 port map( IN1 => n156, IN2 => n157, IN3 => n142, QN => n133);
   U47 : NAND3X1 port map( IN1 => n81, IN2 => n264, IN3 => n75, QN => n94);
   U48 : NBUFFX2 port map( INP => n44, Z => n13);
   U49 : INVX0 port map( INP => cyc_s_1_port, ZN => n14);
   U50 : AND4X1 port map( IN1 => n157, IN2 => n11, IN3 => n81, IN4 => n6, Q => 
                           n15);
   U51 : AND4X1 port map( IN1 => n157, IN2 => n11, IN3 => n81, IN4 => n6, Q => 
                           n16);
   U52 : AO22X2 port map( IN1 => perm_output_60_port, IN2 => n218, IN3 => 
                           cyc_state_update_60_port, IN4 => n50, Q => 
                           ramainput_60_port);
   U53 : AO22X2 port map( IN1 => perm_output_40_port, IN2 => n215, IN3 => 
                           cyc_state_update_40_port, IN4 => n56, Q => 
                           ramainput_40_port);
   U54 : AO22X2 port map( IN1 => perm_output_82_port, IN2 => n221, IN3 => 
                           cyc_state_update_82_port, IN4 => n48, Q => 
                           ramainput_82_port);
   U55 : AO22X2 port map( IN1 => perm_output_83_port, IN2 => n221, IN3 => 
                           cyc_state_update_83_port, IN4 => n48, Q => 
                           ramainput_83_port);
   U56 : AO22X2 port map( IN1 => perm_output_10_port, IN2 => n200, IN3 => 
                           cyc_state_update_10_port, IN4 => n60, Q => 
                           ramainput_10_port);
   U57 : AO22X2 port map( IN1 => perm_output_89_port, IN2 => n222, IN3 => 
                           cyc_state_update_89_port, IN4 => n48, Q => 
                           ramainput_89_port);
   U58 : AO22X2 port map( IN1 => perm_output_62_port, IN2 => n218, IN3 => 
                           cyc_state_update_62_port, IN4 => n50, Q => 
                           ramainput_62_port);
   U59 : AO22X2 port map( IN1 => perm_output_117_port, IN2 => n201, IN3 => 
                           cyc_state_update_117_port, IN4 => n60, Q => 
                           ramainput_117_port);
   U60 : AO22X2 port map( IN1 => perm_output_119_port, IN2 => n201, IN3 => 
                           cyc_state_update_119_port, IN4 => n59, Q => 
                           ramainput_119_port);
   U61 : AO22X2 port map( IN1 => perm_output_63_port, IN2 => n218, IN3 => 
                           cyc_state_update_63_port, IN4 => n50, Q => 
                           ramainput_63_port);
   U62 : AO22X2 port map( IN1 => perm_output_65_port, IN2 => n218, IN3 => 
                           cyc_state_update_65_port, IN4 => n50, Q => 
                           ramainput_65_port);
   U63 : AO22X2 port map( IN1 => perm_output_54_port, IN2 => n217, IN3 => 
                           cyc_state_update_54_port, IN4 => n55, Q => 
                           ramainput_54_port);
   U64 : AO22X2 port map( IN1 => perm_output_55_port, IN2 => n217, IN3 => 
                           cyc_state_update_55_port, IN4 => n55, Q => 
                           ramainput_55_port);
   U65 : AO22X2 port map( IN1 => perm_output_12_port, IN2 => n202, IN3 => 
                           cyc_state_update_12_port, IN4 => n59, Q => 
                           ramainput_12_port);
   U66 : AO22X2 port map( IN1 => perm_output_58_port, IN2 => n217, IN3 => 
                           cyc_state_update_58_port, IN4 => n50, Q => 
                           ramainput_58_port);
   U67 : AO22X2 port map( IN1 => perm_output_106_port, IN2 => n200, IN3 => 
                           cyc_state_update_106_port, IN4 => n61, Q => 
                           ramainput_106_port);
   U68 : AO22X2 port map( IN1 => perm_output_64_port, IN2 => n218, IN3 => 
                           cyc_state_update_64_port, IN4 => n50, Q => 
                           ramainput_64_port);
   U69 : AO22X2 port map( IN1 => perm_output_72_port, IN2 => n220, IN3 => 
                           cyc_state_update_72_port, IN4 => n49, Q => 
                           ramainput_72_port);
   U70 : AO22X2 port map( IN1 => perm_output_42_port, IN2 => n216, IN3 => 
                           cyc_state_update_42_port, IN4 => n56, Q => 
                           ramainput_42_port);
   U71 : AO22X2 port map( IN1 => perm_output_28_port, IN2 => n203, IN3 => 
                           cyc_state_update_28_port, IN4 => n57, Q => 
                           ramainput_28_port);
   U72 : AO22X2 port map( IN1 => perm_output_33_port, IN2 => n214, IN3 => 
                           cyc_state_update_33_port, IN4 => n57, Q => 
                           ramainput_33_port);
   U73 : AO22X2 port map( IN1 => perm_output_74_port, IN2 => n220, IN3 => 
                           cyc_state_update_74_port, IN4 => n49, Q => 
                           ramainput_74_port);
   U74 : AO22X2 port map( IN1 => perm_output_80_port, IN2 => n221, IN3 => 
                           cyc_state_update_80_port, IN4 => n48, Q => 
                           ramainput_80_port);
   U75 : AO22X2 port map( IN1 => perm_output_16_port, IN2 => n202, IN3 => 
                           cyc_state_update_16_port, IN4 => n58, Q => 
                           ramainput_16_port);
   U76 : AO22X2 port map( IN1 => perm_output_19_port, IN2 => n202, IN3 => 
                           cyc_state_update_19_port, IN4 => n58, Q => 
                           ramainput_19_port);
   U77 : AO22X2 port map( IN1 => perm_output_47_port, IN2 => n223, IN3 => 
                           cyc_state_update_47_port, IN4 => n55, Q => 
                           ramainput_47_port);
   U78 : AO22X2 port map( IN1 => perm_output_9_port, IN2 => n62, IN3 => 
                           cyc_state_update_9_port, IN4 => n47, Q => 
                           ramainput_9_port);
   U79 : AO22X2 port map( IN1 => perm_output_110_port, IN2 => n200, IN3 => 
                           cyc_state_update_110_port, IN4 => n60, Q => 
                           ramainput_110_port);
   U80 : AO22X2 port map( IN1 => perm_output_100_port, IN2 => n63, IN3 => 
                           cyc_state_update_100_port, IN4 => n61, Q => 
                           ramainput_100_port);
   U81 : AO22X2 port map( IN1 => perm_output_111_port, IN2 => n200, IN3 => 
                           cyc_state_update_111_port, IN4 => n60, Q => 
                           ramainput_111_port);
   U82 : AO22X2 port map( IN1 => perm_output_114_port, IN2 => n201, IN3 => 
                           cyc_state_update_114_port, IN4 => n60, Q => 
                           ramainput_114_port);
   U83 : AO22X2 port map( IN1 => perm_output_109_port, IN2 => n200, IN3 => 
                           cyc_state_update_109_port, IN4 => n60, Q => 
                           ramainput_109_port);
   U84 : AO22X2 port map( IN1 => perm_output_118_port, IN2 => n201, IN3 => 
                           cyc_state_update_118_port, IN4 => n59, Q => 
                           ramainput_118_port);
   U85 : AO22X2 port map( IN1 => perm_output_56_port, IN2 => n217, IN3 => 
                           cyc_state_update_56_port, IN4 => n55, Q => 
                           ramainput_56_port);
   U86 : AO22X2 port map( IN1 => perm_output_11_port, IN2 => n200, IN3 => 
                           cyc_state_update_11_port, IN4 => n59, Q => 
                           ramainput_11_port);
   U87 : AO22X2 port map( IN1 => perm_output_1_port, IN2 => n202, IN3 => 
                           cyc_state_update_1_port, IN4 => n58, Q => 
                           ramainput_1_port);
   U88 : AO22X2 port map( IN1 => perm_output_23_port, IN2 => n203, IN3 => 
                           cyc_state_update_23_port, IN4 => n58, Q => 
                           ramainput_23_port);
   U89 : AO22X2 port map( IN1 => perm_output_96_port, IN2 => n223, IN3 => 
                           cyc_state_update_96_port, IN4 => n47, Q => 
                           ramainput_96_port);
   U90 : AO22X2 port map( IN1 => perm_output_49_port, IN2 => n217, IN3 => 
                           cyc_state_update_49_port, IN4 => n55, Q => 
                           ramainput_49_port);
   U91 : AO22X2 port map( IN1 => perm_output_14_port, IN2 => n222, IN3 => 
                           cyc_state_update_14_port, IN4 => n58, Q => 
                           ramainput_14_port);
   U92 : AO22X2 port map( IN1 => perm_output_44_port, IN2 => n216, IN3 => 
                           cyc_state_update_44_port, IN4 => n56, Q => 
                           ramainput_44_port);
   U93 : AO22X2 port map( IN1 => perm_output_34_port, IN2 => n214, IN3 => 
                           cyc_state_update_34_port, IN4 => n57, Q => 
                           ramainput_34_port);
   U94 : AO22X2 port map( IN1 => perm_output_46_port, IN2 => n216, IN3 => 
                           cyc_state_update_46_port, IN4 => n55, Q => 
                           ramainput_46_port);
   U95 : AO22X2 port map( IN1 => perm_output_36_port, IN2 => n215, IN3 => 
                           cyc_state_update_36_port, IN4 => n56, Q => 
                           ramainput_36_port);
   U96 : AO22X2 port map( IN1 => perm_output_116_port, IN2 => n201, IN3 => 
                           cyc_state_update_116_port, IN4 => n60, Q => 
                           ramainput_116_port);
   U97 : AO22X2 port map( IN1 => perm_output_17_port, IN2 => n202, IN3 => 
                           cyc_state_update_17_port, IN4 => n58, Q => 
                           ramainput_17_port);
   U98 : AO22X2 port map( IN1 => perm_output_4_port, IN2 => n218, IN3 => 
                           cyc_state_update_4_port, IN4 => n55, Q => 
                           ramainput_4_port);
   U99 : AO22X2 port map( IN1 => perm_output_97_port, IN2 => n223, IN3 => 
                           cyc_state_update_97_port, IN4 => n47, Q => 
                           ramainput_97_port);
   U100 : AO22X2 port map( IN1 => perm_output_105_port, IN2 => n197, IN3 => 
                           cyc_state_update_105_port, IN4 => n61, Q => 
                           ramainput_105_port);
   U101 : DELLN2X2 port map( INP => n147, Z => n17);
   U102 : AO22X2 port map( IN1 => perm_output_86_port, IN2 => n222, IN3 => 
                           cyc_state_update_86_port, IN4 => n48, Q => 
                           ramainput_86_port);
   U103 : AO22X2 port map( IN1 => perm_output_15_port, IN2 => n216, IN3 => 
                           cyc_state_update_15_port, IN4 => n58, Q => 
                           ramainput_15_port);
   U104 : AO22X2 port map( IN1 => perm_output_45_port, IN2 => n216, IN3 => 
                           cyc_state_update_45_port, IN4 => n56, Q => 
                           ramainput_45_port);
   U105 : AO22X2 port map( IN1 => perm_output_18_port, IN2 => n202, IN3 => 
                           cyc_state_update_18_port, IN4 => n58, Q => 
                           ramainput_18_port);
   U106 : AO22X2 port map( IN1 => perm_output_38_port, IN2 => n215, IN3 => 
                           cyc_state_update_38_port, IN4 => n56, Q => 
                           ramainput_38_port);
   U107 : AO22X2 port map( IN1 => perm_output_50_port, IN2 => n219, IN3 => 
                           cyc_state_update_50_port, IN4 => n55, Q => 
                           ramainput_50_port);
   U108 : AO22X2 port map( IN1 => perm_output_73_port, IN2 => n220, IN3 => 
                           cyc_state_update_73_port, IN4 => n49, Q => 
                           ramainput_73_port);
   U109 : AO22X2 port map( IN1 => perm_output_115_port, IN2 => n201, IN3 => 
                           cyc_state_update_115_port, IN4 => n60, Q => 
                           ramainput_115_port);
   U110 : AO22X2 port map( IN1 => perm_output_112_port, IN2 => n201, IN3 => 
                           cyc_state_update_112_port, IN4 => n60, Q => 
                           ramainput_112_port);
   U111 : AO22X2 port map( IN1 => perm_output_79_port, IN2 => n221, IN3 => 
                           cyc_state_update_79_port, IN4 => n48, Q => 
                           ramainput_79_port);
   U112 : AO22X2 port map( IN1 => perm_output_78_port, IN2 => n220, IN3 => 
                           cyc_state_update_78_port, IN4 => n49, Q => 
                           ramainput_78_port);
   U113 : AO22X2 port map( IN1 => perm_output_51_port, IN2 => n216, IN3 => 
                           cyc_state_update_51_port, IN4 => n55, Q => 
                           ramainput_51_port);
   U114 : AO22X2 port map( IN1 => perm_output_61_port, IN2 => n218, IN3 => 
                           cyc_state_update_61_port, IN4 => n50, Q => 
                           ramainput_61_port);
   U115 : AO22X2 port map( IN1 => perm_output_13_port, IN2 => n220, IN3 => 
                           cyc_state_update_13_port, IN4 => n58, Q => 
                           ramainput_13_port);
   U116 : AO22X2 port map( IN1 => perm_output_0_port, IN2 => n216, IN3 => 
                           cyc_state_update_0_port, IN4 => n61, Q => 
                           ramainput_0_port);
   U117 : AO22X2 port map( IN1 => perm_output_53_port, IN2 => n217, IN3 => 
                           cyc_state_update_53_port, IN4 => n55, Q => 
                           ramainput_53_port);
   U118 : AO22X2 port map( IN1 => perm_output_21_port, IN2 => n202, IN3 => 
                           cyc_state_update_21_port, IN4 => n58, Q => 
                           ramainput_21_port);
   U119 : AO22X2 port map( IN1 => perm_output_32_port, IN2 => n214, IN3 => 
                           cyc_state_update_32_port, IN4 => n57, Q => 
                           ramainput_32_port);
   U120 : AO22X2 port map( IN1 => perm_output_59_port, IN2 => n217, IN3 => 
                           cyc_state_update_59_port, IN4 => n50, Q => 
                           ramainput_59_port);
   U121 : AO22X2 port map( IN1 => perm_output_8_port, IN2 => n222, IN3 => 
                           cyc_state_update_8_port, IN4 => n47, Q => 
                           ramainput_8_port);
   U122 : AO22X2 port map( IN1 => perm_output_104_port, IN2 => n197, IN3 => 
                           cyc_state_update_104_port, IN4 => n61, Q => 
                           ramainput_104_port);
   U125 : AO22X2 port map( IN1 => perm_addr_0_port, IN2 => n16, IN3 => n198, 
                           IN4 => dcount_2_port, Q => addrmux2_0_port);
   U126 : NAND3X1 port map( IN1 => n46, IN2 => n13, IN3 => cyc_s_1_port, QN => 
                           n68);
   U127 : NAND2X0 port map( IN1 => n21, IN2 => N275, QN => n18);
   U128 : AND2X1 port map( IN1 => n18, IN2 => n19, Q => N307);
   U129 : OR2X1 port map( IN1 => n20, IN2 => n26, Q => n19);
   U130 : INVX0 port map( INP => n29, ZN => n20);
   U131 : AND2X1 port map( IN1 => n5, IN2 => n29, Q => n21);
   U132 : DELLN2X2 port map( INP => n270, Z => bdo_3_port);
   U133 : DELLN2X2 port map( INP => n271, Z => bdo_1_port);
   U134 : DELLN2X2 port map( INP => n266, Z => bdo_30_port);
   U135 : AO22X2 port map( IN1 => perm_output_84_port, IN2 => n221, IN3 => 
                           cyc_state_update_84_port, IN4 => n48, Q => 
                           ramainput_84_port);
   U136 : DELLN2X2 port map( INP => n269, Z => bdo_5_port);
   U137 : NAND3X4 port map( IN1 => n251, IN2 => n162, IN3 => n231, QN => n160);
   U138 : AND2X4 port map( IN1 => n3, IN2 => n105, Q => n158);
   U139 : AO22X2 port map( IN1 => perm_output_7_port, IN2 => n221, IN3 => 
                           cyc_state_update_7_port, IN4 => n48, Q => 
                           ramainput_7_port);
   U140 : AO22X2 port map( IN1 => perm_output_39_port, IN2 => n215, IN3 => 
                           cyc_state_update_39_port, IN4 => n56, Q => 
                           ramainput_39_port);
   U141 : AO22X2 port map( IN1 => perm_output_71_port, IN2 => n219, IN3 => 
                           cyc_state_update_71_port, IN4 => n49, Q => 
                           ramainput_71_port);
   U142 : AO22X2 port map( IN1 => perm_output_95_port, IN2 => n223, IN3 => 
                           cyc_state_update_95_port, IN4 => n47, Q => 
                           ramainput_95_port);
   U143 : AO22X2 port map( IN1 => perm_output_126_port, IN2 => n214, IN3 => 
                           cyc_state_update_126_port, IN4 => n59, Q => 
                           ramainput_126_port);
   U144 : AO22X2 port map( IN1 => perm_output_35_port, IN2 => n215, IN3 => 
                           cyc_state_update_35_port, IN4 => n56, Q => 
                           ramainput_35_port);
   U145 : AO22X2 port map( IN1 => perm_output_70_port, IN2 => n219, IN3 => 
                           cyc_state_update_70_port, IN4 => n49, Q => 
                           ramainput_70_port);
   U146 : AO22X2 port map( IN1 => perm_output_87_port, IN2 => n222, IN3 => 
                           cyc_state_update_87_port, IN4 => n48, Q => 
                           ramainput_87_port);
   U147 : AO22X2 port map( IN1 => perm_output_69_port, IN2 => n219, IN3 => 
                           cyc_state_update_69_port, IN4 => n49, Q => 
                           ramainput_69_port);
   U148 : AO22X2 port map( IN1 => perm_output_90_port, IN2 => n222, IN3 => 
                           cyc_state_update_90_port, IN4 => n47, Q => 
                           ramainput_90_port);
   U149 : AO22X2 port map( IN1 => perm_output_25_port, IN2 => n203, IN3 => 
                           cyc_state_update_25_port, IN4 => n57, Q => 
                           ramainput_25_port);
   U150 : AO22X2 port map( IN1 => perm_output_2_port, IN2 => n214, IN3 => 
                           cyc_state_update_2_port, IN4 => n57, Q => 
                           ramainput_2_port);
   U151 : AO22X2 port map( IN1 => perm_output_31_port, IN2 => n214, IN3 => 
                           cyc_state_update_31_port, IN4 => n57, Q => 
                           ramainput_31_port);
   U152 : AO22X2 port map( IN1 => perm_output_88_port, IN2 => n222, IN3 => 
                           cyc_state_update_88_port, IN4 => n48, Q => 
                           ramainput_88_port);
   U153 : AO22X2 port map( IN1 => perm_output_30_port, IN2 => n214, IN3 => 
                           cyc_state_update_30_port, IN4 => n57, Q => 
                           ramainput_30_port);
   U154 : AO22X2 port map( IN1 => perm_output_29_port, IN2 => n214, IN3 => 
                           cyc_state_update_29_port, IN4 => n57, Q => 
                           ramainput_29_port);
   U155 : AO22X2 port map( IN1 => perm_output_26_port, IN2 => n203, IN3 => 
                           cyc_state_update_26_port, IN4 => n57, Q => 
                           ramainput_26_port);
   U156 : AO22X2 port map( IN1 => perm_output_57_port, IN2 => n217, IN3 => 
                           cyc_state_update_57_port, IN4 => n50, Q => 
                           ramainput_57_port);
   U157 : NOR2X0 port map( IN1 => n157, IN2 => rst, QN => n26);
   U158 : DELLN2X2 port map( INP => n267, Z => bdo_7_port);
   U159 : AO22X2 port map( IN1 => perm_output_121_port, IN2 => n200, IN3 => 
                           cyc_state_update_121_port, IN4 => n59, Q => 
                           ramainput_121_port);
   U160 : AO22X2 port map( IN1 => perm_output_125_port, IN2 => n215, IN3 => 
                           cyc_state_update_125_port, IN4 => n59, Q => 
                           ramainput_125_port);
   U161 : AO22X2 port map( IN1 => perm_output_20_port, IN2 => n202, IN3 => 
                           cyc_state_update_20_port, IN4 => n58, Q => 
                           ramainput_20_port);
   U162 : DELLN2X2 port map( INP => n268, Z => bdo_6_port);
   U163 : AO22X2 port map( IN1 => perm_output_108_port, IN2 => n200, IN3 => 
                           cyc_state_update_108_port, IN4 => n60, Q => 
                           ramainput_108_port);
   U164 : AO22X2 port map( IN1 => perm_output_77_port, IN2 => n220, IN3 => 
                           cyc_state_update_77_port, IN4 => n49, Q => 
                           ramainput_77_port);
   U165 : AO22X2 port map( IN1 => perm_output_91_port, IN2 => n223, IN3 => 
                           cyc_state_update_91_port, IN4 => n47, Q => 
                           ramainput_91_port);
   U166 : AO22X2 port map( IN1 => perm_output_120_port, IN2 => n201, IN3 => 
                           cyc_state_update_120_port, IN4 => n59, Q => 
                           ramainput_120_port);
   U167 : NAND2X1 port map( IN1 => n264, IN2 => n30, QN => n29);
   U168 : AO22X2 port map( IN1 => perm_output_123_port, IN2 => n201, IN3 => 
                           cyc_state_update_123_port, IN4 => n59, Q => 
                           ramainput_123_port);
   U169 : AO22X2 port map( IN1 => perm_output_67_port, IN2 => n219, IN3 => 
                           cyc_state_update_67_port, IN4 => n50, Q => 
                           ramainput_67_port);
   U170 : AO22X2 port map( IN1 => perm_output_94_port, IN2 => n223, IN3 => 
                           cyc_state_update_94_port, IN4 => n47, Q => 
                           ramainput_94_port);
   U171 : AO22X2 port map( IN1 => perm_output_92_port, IN2 => n223, IN3 => 
                           cyc_state_update_92_port, IN4 => n47, Q => 
                           ramainput_92_port);
   U172 : AO22X2 port map( IN1 => perm_output_81_port, IN2 => n221, IN3 => 
                           cyc_state_update_81_port, IN4 => n48, Q => 
                           ramainput_81_port);
   U173 : AO22X2 port map( IN1 => perm_output_68_port, IN2 => n219, IN3 => 
                           cyc_state_update_68_port, IN4 => n49, Q => 
                           ramainput_68_port);
   U174 : AO22X2 port map( IN1 => perm_output_66_port, IN2 => n219, IN3 => 
                           cyc_state_update_66_port, IN4 => n50, Q => 
                           ramainput_66_port);
   U175 : AO22X2 port map( IN1 => perm_output_6_port, IN2 => n219, IN3 => 
                           cyc_state_update_6_port, IN4 => n49, Q => 
                           ramainput_6_port);
   U176 : AO22X2 port map( IN1 => perm_output_27_port, IN2 => n203, IN3 => 
                           cyc_state_update_27_port, IN4 => n57, Q => 
                           ramainput_27_port);
   U178 : AO22X2 port map( IN1 => perm_output_122_port, IN2 => n215, IN3 => 
                           cyc_state_update_122_port, IN4 => n59, Q => 
                           ramainput_122_port);
   U179 : AO22X2 port map( IN1 => perm_output_127_port, IN2 => n217, IN3 => 
                           cyc_state_update_127_port, IN4 => n59, Q => 
                           ramainput_127_port);
   U180 : AO22X2 port map( IN1 => perm_output_85_port, IN2 => n222, IN3 => 
                           cyc_state_update_85_port, IN4 => n48, Q => 
                           ramainput_85_port);
   U181 : AO22X2 port map( IN1 => perm_output_75_port, IN2 => n220, IN3 => 
                           cyc_state_update_75_port, IN4 => n49, Q => 
                           ramainput_75_port);
   U182 : AO22X2 port map( IN1 => perm_output_98_port, IN2 => n221, IN3 => 
                           cyc_state_update_98_port, IN4 => n47, Q => 
                           ramainput_98_port);
   U183 : AO22X2 port map( IN1 => perm_output_93_port, IN2 => n223, IN3 => 
                           cyc_state_update_93_port, IN4 => n47, Q => 
                           ramainput_93_port);
   U184 : NAND2X1 port map( IN1 => n39, IN2 => n42, QN => n30);
   U185 : IBUFFX16 port map( INP => n10, ZN => n246);
   U186 : DELLN2X2 port map( INP => n265, Z => bdo_31_port);
   U187 : NAND2X0 port map( IN1 => n33, IN2 => n34, QN => n32);
   U188 : IBUFFX16 port map( INP => n32, ZN => n86);
   U189 : AND2X2 port map( IN1 => n44, IN2 => n45, Q => n147);
   U190 : NAND2X0 port map( IN1 => cyc_s_0_port, IN2 => n147, QN => n35);
   U191 : AND3X1 port map( IN1 => cyc_s_0_port, IN2 => n13, IN3 => cyc_s_1_port
                           , Q => n36);
   U192 : NAND2X0 port map( IN1 => bdo_type_3_port, IN2 => bdo_ready, QN => 
                           n171);
   U193 : INVX0 port map( INP => n246, ZN => key_ready_port);
   U195 : INVX0 port map( INP => n63, ZN => n50);
   U196 : INVX0 port map( INP => n63, ZN => n57);
   U197 : INVX0 port map( INP => n197, ZN => n48);
   U198 : INVX0 port map( INP => n63, ZN => n58);
   U199 : INVX0 port map( INP => n197, ZN => n47);
   U200 : INVX0 port map( INP => n63, ZN => n55);
   U201 : INVX0 port map( INP => n63, ZN => n49);
   U202 : INVX0 port map( INP => n63, ZN => n56);
   U203 : INVX0 port map( INP => n178, ZN => bdo_type_0_port);
   U204 : INVX0 port map( INP => n62, ZN => n59);
   U205 : INVX0 port map( INP => n62, ZN => n60);
   U206 : INVX0 port map( INP => n226, ZN => n63);
   U207 : INVX0 port map( INP => n226, ZN => n197);
   U208 : INVX0 port map( INP => n37, ZN => n247);
   U209 : NAND2X0 port map( IN1 => n184, IN2 => n261, QN => n168);
   U210 : INVX0 port map( INP => n62, ZN => n61);
   U211 : INVX0 port map( INP => n225, ZN => n215);
   U212 : INVX0 port map( INP => n225, ZN => n220);
   U213 : INVX0 port map( INP => n224, ZN => n222);
   U214 : INVX0 port map( INP => n224, ZN => n219);
   U215 : INVX0 port map( INP => n224, ZN => n218);
   U216 : INVX0 port map( INP => n224, ZN => n217);
   U217 : INVX0 port map( INP => n226, ZN => n201);
   U218 : INVX0 port map( INP => n224, ZN => n223);
   U219 : INVX0 port map( INP => n225, ZN => n221);
   U220 : INVX0 port map( INP => n225, ZN => n203);
   U221 : INVX0 port map( INP => n225, ZN => n214);
   U222 : INVX0 port map( INP => n226, ZN => n200);
   U223 : INVX0 port map( INP => n225, ZN => n202);
   U224 : INVX0 port map( INP => n224, ZN => n216);
   U225 : INVX0 port map( INP => bdi_size(0), ZN => n241);
   U226 : NAND2X0 port map( IN1 => n158, IN2 => n91, QN => load_rnd);
   U227 : INVX0 port map( INP => bdi_type(0), ZN => n261);
   U228 : INVX0 port map( INP => en_rnd, ZN => n236);
   U229 : INVX0 port map( INP => bdi_size(1), ZN => n239);
   U230 : NOR2X0 port map( IN1 => n111, IN2 => n259, QN => n165);
   U231 : NOR2X0 port map( IN1 => n252, IN2 => n128, QN => n108);
   U232 : INVX0 port map( INP => n225, ZN => n62);
   U233 : INVX0 port map( INP => en_ins, ZN => n226);
   U234 : INVX0 port map( INP => n80, ZN => n245);
   U235 : INVX0 port map( INP => en_ins, ZN => n224);
   U236 : INVX0 port map( INP => en_ins, ZN => n225);
   U237 : INVX0 port map( INP => n83, ZN => n231);
   U238 : INVX0 port map( INP => n84, ZN => n244);
   U239 : INVX0 port map( INP => n94, ZN => n248);
   U240 : INVX0 port map( INP => n149, ZN => n243);
   U241 : NOR2X0 port map( IN1 => dcount_start_value_3, IN2 => n252, QN => n161
                           );
   U242 : NAND2X0 port map( IN1 => n132, IN2 => n251, QN => n174);
   U243 : NAND2X0 port map( IN1 => n251, IN2 => n32, QN => n172);
   U244 : NOR2X0 port map( IN1 => n97, IN2 => n162, QN => n132);
   U245 : INVX0 port map( INP => cu_cd_s_6_port, ZN => n257);
   U246 : NOR2X0 port map( IN1 => n138, IN2 => n142, QN => en_rnd);
   U247 : INVX0 port map( INP => n118, ZN => n259);
   U248 : NAND2X0 port map( IN1 => n264, IN2 => n88, QN => n80);
   U249 : NAND2X0 port map( IN1 => n254, IN2 => n91, QN => n89);
   U250 : NOR2X0 port map( IN1 => n105, IN2 => n137, QN => n128);
   U251 : AND2X1 port map( IN1 => bdi_valid, IN2 => n185, Q => n129);
   U252 : OR2X1 port map( IN1 => n73_port, IN2 => n81, Q => n91);
   U253 : OR2X1 port map( IN1 => n68, IN2 => n185, Q => n111);
   U254 : NAND2X0 port map( IN1 => n80, IN2 => n82, QN => n76);
   U256 : NAND2X0 port map( IN1 => n84, IN2 => n162, QN => n96);
   U259 : NAND2X0 port map( IN1 => n142, IN2 => n96, QN => en_ins);
   U279 : NAND2X0 port map( IN1 => n163, IN2 => n232, QN => n83);
   U281 : NAND2X1 port map( IN1 => n249, IN2 => n115, QN => n113);
   U294 : INVX0 port map( INP => n90, ZN => n252);
   U295 : INVX0 port map( INP => n68, ZN => n250);
   U298 : NAND2X0 port map( IN1 => msg_auth_ready, IN2 => bdi_valid, QN => n149
                           );
   U299 : INVX0 port map( INP => n142, ZN => n249);
   U311 : NAND2X0 port map( IN1 => n264, IN2 => n154, QN => n150);
   U322 : NAND4X0 port map( IN1 => n90, IN2 => n37, IN3 => n81, IN4 => n155, QN
                           => n154);
   U325 : NOR2X0 port map( IN1 => n250, IN2 => n133, QN => n155);
   U327 : INVX0 port map( INP => n140, ZN => n233);
   U332 : AND2X1 port map( IN1 => n69, IN2 => n68, Q => n39);
   U336 : NOR4X0 port map( IN1 => n258, IN2 => n115, IN3 => n138, IN4 => n142, 
                           QN => ins_start_value_0);
   U345 : INVX0 port map( INP => n104, ZN => n258);
   U347 : NAND2X0 port map( IN1 => n148, IN2 => cyc_s_0_port, QN => n157);
   U348 : INVX0 port map( INP => n66, ZN => n255);
   U349 : NAND2X0 port map( IN1 => n65, IN2 => n3, QN => cu_cd_s_1);
   U350 : INVX0 port map( INP => n65, ZN => n253);
   U351 : NOR2X0 port map( IN1 => n232, IN2 => n235, QN => n176);
   U352 : INVX0 port map( INP => dcount_0_port, ZN => n232);
   U354 : NAND2X0 port map( IN1 => n148, IN2 => n46, QN => n142);
   U355 : INVX0 port map( INP => bdi_type(1), ZN => n263);
   U356 : AND4X1 port map( IN1 => bdi_valid, IN2 => n187, IN3 => n73_port, IN4 
                           => n240, Q => n186);
   U357 : INVX0 port map( INP => n188, ZN => n240);
   U359 : INVX0 port map( INP => dcount_3_port, ZN => n235);
   U360 : NAND3X0 port map( IN1 => calling_state_0_port, IN2 => n51, IN3 => 
                           calling_state_1_port, QN => n137);
   U361 : INVX0 port map( INP => dcount_2_port, ZN => n234);
   U365 : NAND3X0 port map( IN1 => n52, IN2 => n51, IN3 => calling_state_0_port
                           , QN => n118);
   U366 : NAND2X0 port map( IN1 => n78, IN2 => n79, QN => n206);
   U367 : NAND3X0 port map( IN1 => n80, IN2 => n260, IN3 => n72_port, QN => n79
                           );
   U368 : NAND2X0 port map( IN1 => en_rnd, IN2 => n115, QN => n135);
   U369 : NOR2X0 port map( IN1 => n259, IN2 => n245, QN => n77);
   U370 : NOR2X0 port map( IN1 => n157, IN2 => decrypt_op_s, QN => 
                           bdo_type_3_port);
   U371 : NOR2X0 port map( IN1 => n231, IN2 => n51, QN => n87);
   U372 : INVX0 port map( INP => rnd_counter_2_port, ZN => n237);
   U373 : NOR2X0 port map( IN1 => n98, IN2 => rst, QN => n99);
   U374 : NOR2X0 port map( IN1 => n164, IN2 => n140, QN => end_of_block);
   U375 : NOR2X0 port map( IN1 => n157, IN2 => n54, QN => n141);
   U376 : NOR2X0 port map( IN1 => n94, IN2 => n90, QN => n93);
   U377 : NOR2X0 port map( IN1 => dcount_2_port, IN2 => dcount_0_port, QN => 
                           n122);
   U378 : NAND2X0 port map( IN1 => dcount_0_port, IN2 => n163, QN => n140);
   U379 : AO22X1 port map( IN1 => n71, IN2 => gtr_one_perm, IN3 => n72_port, 
                           IN4 => n73_port, Q => n204);
   U380 : AOI21X1 port map( IN1 => n41, IN2 => n75, IN3 => rst, QN => n71);
   U381 : INVX0 port map( INP => rst, ZN => n264);
   U382 : NOR2X0 port map( IN1 => n81, IN2 => rst, QN => n72_port);
   U383 : NBUFFX2 port map( INP => clk, Z => n40);
   U384 : NOR2X0 port map( IN1 => bdi_size(1), IN2 => bdi_size(0), QN => n188);
   U385 : NOR2X0 port map( IN1 => n167, IN2 => n168, QN => n166);
   U386 : NAND2X0 port map( IN1 => n170, IN2 => n167, QN => bdi_ready);
   U387 : NAND2X0 port map( IN1 => n36, IN2 => n186, QN => n167);
   U388 : NAND2X0 port map( IN1 => key_update_internal_0_port, IN2 => n31, QN 
                           => n162);
   U389 : INVX0 port map( INP => n2, ZN => n41);
   U390 : INVX0 port map( INP => n70, ZN => n238);
   U391 : NOR3X0 port map( IN1 => bdo_type_3_port, IN2 => n254, IN3 => n256, QN
                           => n42);
   U392 : INVX0 port map( INP => n156, ZN => n256);
   U393 : INVX0 port map( INP => n81, ZN => n254);
   U394 : INVX0 port map( INP => bdi_type(2), ZN => n262);
   U395 : NAND3X1 port map( IN1 => n46, IN2 => n14, IN3 => cyc_s_2_port, QN => 
                           n81);
   U396 : NAND3X1 port map( IN1 => cyc_s_0_port, IN2 => cyc_s_2_port, IN3 => 
                           n45, QN => n156);
   U397 : NAND2X0 port map( IN1 => bdo_ready, IN2 => n242, QN => n124);
   U398 : NAND2X1 port map( IN1 => n178, IN2 => n179, QN => 
                           cyc_state_update_sel_1_port);
   U399 : NAND2X0 port map( IN1 => n183, IN2 => n168, QN => n178);
   U400 : NOR2X0 port map( IN1 => n260, IN2 => calling_state_1_port, QN => n185
                           );
   U401 : NOR2X0 port map( IN1 => n52, IN2 => n260, QN => n189);
   U402 : NOR2X0 port map( IN1 => n83, IN2 => n86, QN => n152);
   U403 : INVX0 port map( INP => n180, ZN => n260);
   U404 : NOR2X0 port map( IN1 => key_valid, IN2 => bdi_valid, QN => n146);
   U405 : NAND2X0 port map( IN1 => key_valid, IN2 => N103, QN => n175);
   U406 : NOR2X0 port map( IN1 => key_valid, IN2 => bdi_eot, QN => n121);
   U407 : INVX0 port map( INP => n121, ZN => n242);
   U408 : NAND2X0 port map( IN1 => n146, IN2 => n17, QN => n145);
   U409 : NOR2X0 port map( IN1 => n41, IN2 => n86, QN => n84);
   U410 : NOR2X0 port map( IN1 => calling_state_2_port, IN2 => 
                           calling_state_0_port, QN => n180);
   U411 : NOR2X0 port map( IN1 => n177, IN2 => n239, QN => cycd_sel_1_port);
   U412 : NAND2X0 port map( IN1 => cyc_s_0_port, IN2 => n147, QN => n74);
   U413 : NAND2X0 port map( IN1 => n17, IN2 => n46, QN => n90);
   U414 : NOR2X0 port map( IN1 => n250, IN2 => n230, QN => n177);
   U415 : INVX0 port map( INP => n167, ZN => n230);
   U416 : NOR2X0 port map( IN1 => n177, IN2 => n241, QN => cycd_sel_0_port);
   U417 : NOR2X0 port map( IN1 => addr_sel_1_port, IN2 => n12, QN => n198);
   U418 : NAND2X0 port map( IN1 => key_ready_port, IN2 => n97, QN => n95);
   U419 : AOI21X1 port map( IN1 => dcount_2_port, IN2 => dcount_1_port, IN3 => 
                           dcount_3_port, QN => N73);
   U420 : AO21X1 port map( IN1 => dcount_1_port, IN2 => dcount_0_port, IN3 => 
                           dcount_2_port, Q => n227);
   U421 : NAND2X0 port map( IN1 => dcount_3_port, IN2 => n227, QN => N72);
   U422 : NOR2X0 port map( IN1 => dcount_3_port, IN2 => dcount_2_port, QN => 
                           N103);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_LWC_1.all;

entity PreProcessor_1 is

   port( clk, rst : in std_logic;  pdi_data : in std_logic_vector (31 downto 0)
         ;  pdi_valid : in std_logic;  pdi_ready : out std_logic;  sdi_data : 
         in std_logic_vector (31 downto 0);  sdi_valid : in std_logic;  
         sdi_ready : out std_logic;  key : out std_logic_vector (31 downto 0); 
         key_valid : out std_logic;  key_ready : in std_logic;  bdi : out 
         std_logic_vector (31 downto 0);  bdi_valid : out std_logic;  bdi_ready
         : in std_logic;  bdi_pad_loc, bdi_valid_bytes : out std_logic_vector 
         (3 downto 0);  bdi_size : out std_logic_vector (2 downto 0);  bdi_eot,
         bdi_eoi : out std_logic;  bdi_type : out std_logic_vector (3 downto 0)
         ;  decrypt, hash, key_update : out std_logic;  cmd : out 
         std_logic_vector (31 downto 0);  cmd_valid : out std_logic;  cmd_ready
         : in std_logic);

end PreProcessor_1;

architecture SYN_PreProcessor of PreProcessor_1 is

   component AND4X1
      port( IN1, IN2, IN3, IN4 : in std_logic;  Q : out std_logic);
   end component;
   
   component NOR4X0
      port( IN1, IN2, IN3, IN4 : in std_logic;  QN : out std_logic);
   end component;
   
   component NOR3X0
      port( IN1, IN2, IN3 : in std_logic;  QN : out std_logic);
   end component;
   
   component OA21X1
      port( IN1, IN2, IN3 : in std_logic;  Q : out std_logic);
   end component;
   
   component NAND2X0
      port( IN1, IN2 : in std_logic;  QN : out std_logic);
   end component;
   
   component AND2X2
      port( IN1, IN2 : in std_logic;  Q : out std_logic);
   end component;
   
   component NOR2X0
      port( IN1, IN2 : in std_logic;  QN : out std_logic);
   end component;
   
   component INVX0
      port( INP : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3X0
      port( IN1, IN2, IN3 : in std_logic;  QN : out std_logic);
   end component;
   
   component NAND2X1
      port( IN1, IN2 : in std_logic;  QN : out std_logic);
   end component;
   
   component AND2X1
      port( IN1, IN2 : in std_logic;  Q : out std_logic);
   end component;
   
   component DATA_PISO_1
      port( clk, rst : in std_logic;  data_size_p : in std_logic_vector (2 
            downto 0);  data_size_s : out std_logic_vector (2 downto 0);  
            data_s : out std_logic_vector (31 downto 0);  data_valid_s : out 
            std_logic;  data_ready_s : in std_logic;  data_p : in 
            std_logic_vector (31 downto 0);  data_valid_p : in std_logic;  
            data_ready_p : out std_logic;  valid_bytes_p : in std_logic_vector 
            (3 downto 0);  valid_bytes_s : out std_logic_vector (3 downto 0);  
            pad_loc_p : in std_logic_vector (3 downto 0);  pad_loc_s : out 
            std_logic_vector (3 downto 0);  eoi_p : in std_logic;  eoi_s : out 
            std_logic;  eot_p : in std_logic;  eot_s : out std_logic);
   end component;
   
   component KEY_PISO_1
      port( clk, rst : in std_logic;  data_s : out std_logic_vector (31 downto 
            0);  data_valid_s : out std_logic;  data_ready_s : in std_logic;  
            data_p : in std_logic_vector (31 downto 0);  data_valid_p : in 
            std_logic;  data_ready_p : out std_logic);
   end component;
   
   component StepDownCountLd_N16_step4_1_0
      port( clk, len, ena : in std_logic;  load : in std_logic_vector (15 
            downto 0);  count : out std_logic_vector (15 downto 0));
   end component;
   
   component OR4X1
      port( IN1, IN2, IN3, IN4 : in std_logic;  Q : out std_logic);
   end component;
   
   component OR2X1
      port( IN1, IN2 : in std_logic;  Q : out std_logic);
   end component;
   
   component NAND4X0
      port( IN1, IN2, IN3, IN4 : in std_logic;  QN : out std_logic);
   end component;
   
   component AO222X1
      port( IN1, IN2, IN3, IN4, IN5, IN6 : in std_logic;  Q : out std_logic);
   end component;
   
   component OA22X1
      port( IN1, IN2, IN3, IN4 : in std_logic;  Q : out std_logic);
   end component;
   
   component OAI22X1
      port( IN1, IN2, IN3, IN4 : in std_logic;  QN : out std_logic);
   end component;
   
   component OAI21X1
      port( IN1, IN2, IN3 : in std_logic;  QN : out std_logic);
   end component;
   
   component AO22X1
      port( IN1, IN2, IN3, IN4 : in std_logic;  Q : out std_logic);
   end component;
   
   component AOI221X1
      port( IN1, IN2, IN3, IN4, IN5 : in std_logic;  QN : out std_logic);
   end component;
   
   component AO221X1
      port( IN1, IN2, IN3, IN4, IN5 : in std_logic;  Q : out std_logic);
   end component;
   
   component AO21X1
      port( IN1, IN2, IN3 : in std_logic;  Q : out std_logic);
   end component;
   
   component AND3X1
      port( IN1, IN2, IN3 : in std_logic;  Q : out std_logic);
   end component;
   
   component DFFX1
      port( D, CLK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal bdi_type_3_port, bdi_type_2_port, bdi_type_0_port, decrypt_port, 
      hash_port, key_update_port, len_SegLenCnt, en_SegLenCnt, 
      load_SegLenCnt_15_port, load_SegLenCnt_14_port, load_SegLenCnt_13_port, 
      load_SegLenCnt_12_port, load_SegLenCnt_11_port, load_SegLenCnt_10_port, 
      load_SegLenCnt_9_port, load_SegLenCnt_8_port, load_SegLenCnt_7_port, 
      load_SegLenCnt_6_port, load_SegLenCnt_5_port, load_SegLenCnt_4_port, 
      load_SegLenCnt_3_port, load_SegLenCnt_2_port, load_SegLenCnt_1_port, 
      load_SegLenCnt_0_port, dout_SegLenCnt_15_port, dout_SegLenCnt_14_port, 
      dout_SegLenCnt_13_port, dout_SegLenCnt_12_port, dout_SegLenCnt_11_port, 
      dout_SegLenCnt_10_port, dout_SegLenCnt_9_port, dout_SegLenCnt_8_port, 
      dout_SegLenCnt_7_port, dout_SegLenCnt_6_port, dout_SegLenCnt_5_port, 
      dout_SegLenCnt_4_port, dout_SegLenCnt_3_port, dout_SegLenCnt_2_port, 
      dout_SegLenCnt_1_port, dout_SegLenCnt_0_port, N64, 
      bdi_valid_bytes_p_3_port, bdi_valid_bytes_p_1_port, 
      bdi_valid_bytes_p_0_port, bdi_pad_loc_p_3_port, bdi_pad_loc_p_1_port, 
      bdi_pad_loc_p_0_port, eoi_flag, eot_flag, bdi_size_p_2_port, 
      bdi_size_p_1_port, bdi_size_p_0_port, bdi_eoi_internal, bdi_eot_internal,
      key_ready_p, key_valid_p, bdi_ready_p, bdi_valid_p, pr_state_3_port, 
      pr_state_2_port, pr_state_1_port, pr_state_0_port, N206, N207, N208, N209
      , n12, n27, n28, n29, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, 
      n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61
      , n62, n63, n64_port, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, 
      n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89
      , n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, 
      n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, 
      n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, 
      n127, n128, n129, n130, n131, n132, n1, n2, n3, n4, n5, n6, n7, n8, n9, 
      n10, n11, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, 
      bdi_type_1_port, n25, n26, n30, n31, n32, n33, n34, n35, n36, n133, n134,
      n_3231, n_3232, n_3233, n_3234 : std_logic;

begin
   bdi_type <= ( bdi_type_3_port, bdi_type_2_port, bdi_type_1_port, 
      bdi_type_0_port );
   decrypt <= decrypt_port;
   hash <= hash_port;
   key_update <= key_update_port;
   cmd <= ( pdi_data(31), pdi_data(30), pdi_data(29), pdi_data(28), 
      pdi_data(27), pdi_data(26), pdi_data(25), pdi_data(24), pdi_data(23), 
      pdi_data(22), pdi_data(21), pdi_data(20), pdi_data(19), pdi_data(18), 
      pdi_data(17), pdi_data(16), pdi_data(15), pdi_data(14), pdi_data(13), 
      pdi_data(12), pdi_data(11), pdi_data(10), pdi_data(9), pdi_data(8), 
      pdi_data(7), pdi_data(6), pdi_data(5), pdi_data(4), pdi_data(3), 
      pdi_data(2), pdi_data(1), pdi_data(0) );
   
   pr_state_reg_0_inst : DFFX1 port map( D => N206, CLK => clk, Q => 
                           pr_state_0_port, QN => n29);
   eoi_flag_reg : DFFX1 port map( D => n130, CLK => clk, Q => eoi_flag, QN => 
                           n_3231);
   eot_flag_reg : DFFX1 port map( D => n129, CLK => clk, Q => eot_flag, QN => 
                           n_3232);
   pr_state_reg_1_inst : DFFX1 port map( D => N207, CLK => clk, Q => 
                           pr_state_1_port, QN => n28);
   pr_state_reg_2_inst : DFFX1 port map( D => N208, CLK => clk, Q => 
                           pr_state_2_port, QN => n_3233);
   pr_state_reg_3_inst : DFFX1 port map( D => N209, CLK => clk, Q => 
                           pr_state_3_port, QN => n27);
   decrypt_internal_reg : DFFX1 port map( D => n131, CLK => clk, Q => 
                           decrypt_port, QN => n12);
   hash_internal_reg : DFFX1 port map( D => n132, CLK => clk, Q => hash_port, 
                           QN => n_3234);
   U79 : NAND3X0 port map( IN1 => n1, IN2 => n38, IN3 => n39, QN => sdi_ready);
   U80 : AO221X1 port map( IN1 => bdi_ready_p, IN2 => n40, IN3 => n41, IN4 => 
                           n42, IN5 => n43, Q => pdi_ready);
   U81 : AO21X1 port map( IN1 => cmd_ready, IN2 => n25, IN3 => n44, Q => n43);
   U82 : NAND3X0 port map( IN1 => n45, IN2 => n17, IN3 => pdi_valid, QN => n42)
                           ;
   U83 : OR2X1 port map( IN1 => n46, IN2 => n34, Q => n45);
   U84 : AO22X1 port map( IN1 => pdi_data(25), IN2 => n16, IN3 => eot_flag, IN4
                           => n47, Q => n129);
   U85 : AO22X1 port map( IN1 => pdi_data(26), IN2 => n16, IN3 => eoi_flag, IN4
                           => n47, Q => n130);
   U86 : NAND4X0 port map( IN1 => n37, IN2 => n38, IN3 => n48, IN4 => n49, QN 
                           => n47);
   U87 : NOR3X0 port map( IN1 => n57, IN2 => bdi_type_1_port, IN3 => n41, QN =>
                           n48);
   U88 : AO22X1 port map( IN1 => decrypt_port, IN2 => n20, IN3 => pdi_data(28),
                           IN4 => n58, Q => n131);
   U89 : NOR3X0 port map( IN1 => n59, IN2 => n133, IN3 => n60, QN => n58);
   U90 : AO22X1 port map( IN1 => hash_port, IN2 => n59, IN3 => n61, IN4 => n46,
                           Q => n132);
   U91 : NAND4X0 port map( IN1 => n56, IN2 => n37, IN3 => n26, IN4 => n62, QN 
                           => n59);
   U92 : NOR3X0 port map( IN1 => n23, IN2 => bdi_type_2_port, IN3 => n57, QN =>
                           n62);
   U93 : AO22X1 port map( IN1 => pdi_data(9), IN2 => n1, IN3 => sdi_data(9), 
                           IN4 => n31, Q => load_SegLenCnt_9_port);
   U94 : AO22X1 port map( IN1 => pdi_data(8), IN2 => n37, IN3 => sdi_data(8), 
                           IN4 => n31, Q => load_SegLenCnt_8_port);
   U95 : AO22X1 port map( IN1 => pdi_data(7), IN2 => n1, IN3 => sdi_data(7), 
                           IN4 => n31, Q => load_SegLenCnt_7_port);
   U96 : AO22X1 port map( IN1 => pdi_data(6), IN2 => n37, IN3 => sdi_data(6), 
                           IN4 => n31, Q => load_SegLenCnt_6_port);
   U97 : AO22X1 port map( IN1 => pdi_data(5), IN2 => n1, IN3 => sdi_data(5), 
                           IN4 => n31, Q => load_SegLenCnt_5_port);
   U98 : AO22X1 port map( IN1 => pdi_data(4), IN2 => n37, IN3 => sdi_data(4), 
                           IN4 => n31, Q => load_SegLenCnt_4_port);
   U99 : AO22X1 port map( IN1 => pdi_data(3), IN2 => n1, IN3 => sdi_data(3), 
                           IN4 => n31, Q => load_SegLenCnt_3_port);
   U100 : AO22X1 port map( IN1 => pdi_data(2), IN2 => n37, IN3 => sdi_data(2), 
                           IN4 => n31, Q => load_SegLenCnt_2_port);
   U101 : AO22X1 port map( IN1 => pdi_data(1), IN2 => n1, IN3 => sdi_data(1), 
                           IN4 => n31, Q => load_SegLenCnt_1_port);
   U102 : AO22X1 port map( IN1 => pdi_data(15), IN2 => n37, IN3 => sdi_data(15)
                           , IN4 => n31, Q => load_SegLenCnt_15_port);
   U103 : AO22X1 port map( IN1 => pdi_data(14), IN2 => n1, IN3 => sdi_data(14),
                           IN4 => n31, Q => load_SegLenCnt_14_port);
   U104 : AO22X1 port map( IN1 => pdi_data(13), IN2 => n37, IN3 => sdi_data(13)
                           , IN4 => n31, Q => load_SegLenCnt_13_port);
   U105 : AO22X1 port map( IN1 => pdi_data(12), IN2 => n1, IN3 => sdi_data(12),
                           IN4 => n31, Q => load_SegLenCnt_12_port);
   U106 : AO22X1 port map( IN1 => pdi_data(11), IN2 => n37, IN3 => sdi_data(11)
                           , IN4 => n31, Q => load_SegLenCnt_11_port);
   U107 : AO22X1 port map( IN1 => pdi_data(10), IN2 => n1, IN3 => sdi_data(10),
                           IN4 => n31, Q => load_SegLenCnt_10_port);
   U108 : AO22X1 port map( IN1 => pdi_data(0), IN2 => n1, IN3 => sdi_data(0), 
                           IN4 => n31, Q => load_SegLenCnt_0_port);
   U109 : AO221X1 port map( IN1 => pdi_valid, IN2 => n44, IN3 => sdi_valid, IN4
                           => n31, IN5 => n63, Q => len_SegLenCnt);
   U110 : NAND4X0 port map( IN1 => n64_port, IN2 => n65, IN3 => n66, IN4 => n53
                           , QN => n44);
   U111 : AO22X1 port map( IN1 => key_valid_p, IN2 => key_ready_p, IN3 => n67, 
                           IN4 => pdi_valid, Q => en_SegLenCnt);
   U112 : AND2X1 port map( IN1 => n40, IN2 => bdi_ready_p, Q => n67);
   U114 : OA21X1 port map( IN1 => n68, IN2 => n25, IN3 => pdi_valid, Q => 
                           cmd_valid);
   U115 : OA21X1 port map( IN1 => n46, IN2 => n34, IN3 => n41, Q => n68);
   U116 : AO21X1 port map( IN1 => pdi_valid, IN2 => n40, IN3 => n69, Q => 
                           bdi_valid_p);
   U117 : NAND4X0 port map( IN1 => n70, IN2 => n71, IN3 => n72, IN4 => n73, QN 
                           => n40);
   U118 : OR2X1 port map( IN1 => n12, IN2 => n74, Q => n71);
   U119 : OR2X1 port map( IN1 => bdi_pad_loc_p_0_port, IN2 => 
                           bdi_valid_bytes_p_0_port, Q => 
                           bdi_valid_bytes_p_1_port);
   U120 : NAND3X0 port map( IN1 => n73, IN2 => n77, IN3 => n54, QN => 
                           bdi_type_2_port);
   U121 : NAND4X0 port map( IN1 => n72, IN2 => n73, IN3 => n78, IN4 => n77, QN 
                           => bdi_type_0_port);
   U122 : OR2X1 port map( IN1 => n10, IN2 => dout_SegLenCnt_2_port, Q => 
                           bdi_size_p_2_port);
   U123 : AND3X1 port map( IN1 => n13, IN2 => n15, IN3 => n80, Q => 
                           bdi_pad_loc_p_3_port);
   U124 : NAND3X0 port map( IN1 => n80, IN2 => n15, IN3 => 
                           dout_SegLenCnt_0_port, QN => n75);
   U125 : AND3X1 port map( IN1 => n80, IN2 => n13, IN3 => dout_SegLenCnt_1_port
                           , Q => bdi_pad_loc_p_1_port);
   U126 : AND3X1 port map( IN1 => dout_SegLenCnt_0_port, IN2 => n80, IN3 => 
                           dout_SegLenCnt_1_port, Q => bdi_pad_loc_p_0_port);
   U127 : AND4X1 port map( IN1 => n81, IN2 => n82, IN3 => n83, IN4 => n84, Q =>
                           n80);
   U128 : NOR3X0 port map( IN1 => dout_SegLenCnt_3_port, IN2 => 
                           dout_SegLenCnt_5_port, IN3 => dout_SegLenCnt_4_port,
                           QN => n83);
   U129 : NOR3X0 port map( IN1 => dout_SegLenCnt_10_port, IN2 => 
                           dout_SegLenCnt_12_port, IN3 => 
                           dout_SegLenCnt_11_port, QN => n81);
   U130 : AND2X1 port map( IN1 => eot_flag, IN2 => N64, Q => bdi_eot_internal);
   U131 : AND2X1 port map( IN1 => eoi_flag, IN2 => N64, Q => bdi_eoi_internal);
   U132 : OA21X1 port map( IN1 => n85, IN2 => n86, IN3 => n33, Q => N209);
   U133 : AO221X1 port map( IN1 => n87, IN2 => n21, IN3 => n69, IN4 => n7, IN5 
                           => n88, Q => n86);
   U134 : AO21X1 port map( IN1 => n19, IN2 => n8, IN3 => n89, Q => n88);
   U135 : AO221X1 port map( IN1 => n90, IN2 => n32, IN3 => n25, IN4 => n91, IN5
                           => n92, Q => n85);
   U136 : NAND3X0 port map( IN1 => n64_port, IN2 => n78, IN3 => n93, QN => n92)
                           ;
   U137 : NAND3X0 port map( IN1 => n46, IN2 => n41, IN3 => n55, QN => n93);
   U138 : NAND3X0 port map( IN1 => n55, IN2 => n12, IN3 => n32, QN => n91);
   U139 : AND4X1 port map( IN1 => n95, IN2 => n64_port, IN3 => n73, IN4 => n66,
                           Q => n94);
   U140 : AOI221X1 port map( IN1 => n41, IN2 => n96, IN3 => n79, IN4 => n87, 
                           IN5 => n97, QN => n95);
   U141 : AO22X1 port map( IN1 => n55, IN2 => n34, IN3 => n55, IN4 => n46, Q =>
                           n96);
   U142 : NAND3X0 port map( IN1 => n36, IN2 => n35, IN3 => pdi_data(29), QN => 
                           n60);
   U143 : AO222X1 port map( IN1 => n69, IN2 => n7, IN3 => n30, IN4 => n101, IN5
                           => n19, IN6 => n87, Q => n97);
   U144 : AND2X1 port map( IN1 => n102, IN2 => n103, Q => n69);
   U145 : OAI21X1 port map( IN1 => n74, IN2 => n9, IN3 => n53, QN => n89);
   U146 : OAI22X1 port map( IN1 => n38, IN2 => n134, IN3 => n73, IN4 => n104, 
                           QN => n100);
   U147 : NAND4X0 port map( IN1 => n105, IN2 => n1, IN3 => n106, IN4 => n107, 
                           QN => n99);
   U148 : OA22X1 port map( IN1 => n64_port, IN2 => n108, IN3 => n87, IN4 => n78
                           , Q => n107);
   U150 : NAND3X0 port map( IN1 => n32, IN2 => decrypt_port, IN3 => n63, QN => 
                           n105);
   U151 : OA21X1 port map( IN1 => n112, IN2 => n113, IN3 => n33, Q => N206);
   U152 : AO222X1 port map( IN1 => sdi_valid, IN2 => n31, IN3 => 
                           key_update_port, IN4 => n111, IN5 => n23, IN6 => 
                           n134, Q => n113);
   U154 : AND2X1 port map( IN1 => n57, IN2 => n110, Q => key_update_port);
   U155 : AO222X1 port map( IN1 => n63, IN2 => n115, IN3 => n116, IN4 => n104, 
                           IN5 => pdi_valid, IN6 => n117, Q => n112);
   U156 : NAND4X0 port map( IN1 => n66, IN2 => n53, IN3 => n118, IN4 => n119, 
                           QN => n117);
   U157 : OA21X1 port map( IN1 => n32, IN2 => n65, IN3 => n120, Q => n119);
   U158 : NAND4X0 port map( IN1 => pdi_data(29), IN2 => n35, IN3 => n41, IN4 =>
                           n121, QN => n120);
   U159 : AND2X1 port map( IN1 => pdi_data(28), IN2 => pdi_data(30), Q => n121)
                           ;
   U161 : OR2X1 port map( IN1 => n64_port, IN2 => n109, Q => n118);
   U162 : NAND3X0 port map( IN1 => pdi_valid, IN2 => bdi_ready_p, IN3 => N64, 
                           QN => n104);
   U163 : AND2X1 port map( IN1 => n102, IN2 => n114, Q => n79);
   U164 : AND2X1 port map( IN1 => pr_state_2_port, IN2 => pr_state_3_port, Q =>
                           n102);
   U165 : AND2X1 port map( IN1 => pr_state_2_port, IN2 => n27, Q => n123);
   U166 : OR4X1 port map( IN1 => pdi_data(2), IN2 => pdi_data(3), IN3 => 
                           pdi_data(4), IN4 => pdi_data(5), Q => n128);
   U167 : OR4X1 port map( IN1 => pdi_data(6), IN2 => pdi_data(7), IN3 => 
                           pdi_data(8), IN4 => pdi_data(9), Q => n127);
   U168 : OR4X1 port map( IN1 => pdi_data(0), IN2 => pdi_data(10), IN3 => 
                           pdi_data(11), IN4 => pdi_data(12), Q => n126);
   U169 : OR4X1 port map( IN1 => pdi_data(13), IN2 => pdi_data(14), IN3 => 
                           pdi_data(15), IN4 => pdi_data(1), Q => n125);
   U170 : AND2X1 port map( IN1 => n55, IN2 => n25, Q => n63);
   SegLen : StepDownCountLd_N16_step4_1_0 port map( clk => clk, len => 
                           len_SegLenCnt, ena => en_SegLenCnt, load(15) => 
                           load_SegLenCnt_15_port, load(14) => 
                           load_SegLenCnt_14_port, load(13) => 
                           load_SegLenCnt_13_port, load(12) => 
                           load_SegLenCnt_12_port, load(11) => 
                           load_SegLenCnt_11_port, load(10) => 
                           load_SegLenCnt_10_port, load(9) => 
                           load_SegLenCnt_9_port, load(8) => 
                           load_SegLenCnt_8_port, load(7) => 
                           load_SegLenCnt_7_port, load(6) => 
                           load_SegLenCnt_6_port, load(5) => 
                           load_SegLenCnt_5_port, load(4) => 
                           load_SegLenCnt_4_port, load(3) => 
                           load_SegLenCnt_3_port, load(2) => 
                           load_SegLenCnt_2_port, load(1) => 
                           load_SegLenCnt_1_port, load(0) => 
                           load_SegLenCnt_0_port, count(15) => 
                           dout_SegLenCnt_15_port, count(14) => 
                           dout_SegLenCnt_14_port, count(13) => 
                           dout_SegLenCnt_13_port, count(12) => 
                           dout_SegLenCnt_12_port, count(11) => 
                           dout_SegLenCnt_11_port, count(10) => 
                           dout_SegLenCnt_10_port, count(9) => 
                           dout_SegLenCnt_9_port, count(8) => 
                           dout_SegLenCnt_8_port, count(7) => 
                           dout_SegLenCnt_7_port, count(6) => 
                           dout_SegLenCnt_6_port, count(5) => 
                           dout_SegLenCnt_5_port, count(4) => 
                           dout_SegLenCnt_4_port, count(3) => 
                           dout_SegLenCnt_3_port, count(2) => 
                           dout_SegLenCnt_2_port, count(1) => 
                           dout_SegLenCnt_1_port, count(0) => 
                           dout_SegLenCnt_0_port);
   keyPISO : KEY_PISO_1 port map( clk => clk, rst => rst, data_s(31) => key(31)
                           , data_s(30) => key(30), data_s(29) => key(29), 
                           data_s(28) => key(28), data_s(27) => key(27), 
                           data_s(26) => key(26), data_s(25) => key(25), 
                           data_s(24) => key(24), data_s(23) => key(23), 
                           data_s(22) => key(22), data_s(21) => key(21), 
                           data_s(20) => key(20), data_s(19) => key(19), 
                           data_s(18) => key(18), data_s(17) => key(17), 
                           data_s(16) => key(16), data_s(15) => key(15), 
                           data_s(14) => key(14), data_s(13) => key(13), 
                           data_s(12) => key(12), data_s(11) => key(11), 
                           data_s(10) => key(10), data_s(9) => key(9), 
                           data_s(8) => key(8), data_s(7) => key(7), data_s(6) 
                           => key(6), data_s(5) => key(5), data_s(4) => key(4),
                           data_s(3) => key(3), data_s(2) => key(2), data_s(1) 
                           => key(1), data_s(0) => key(0), data_valid_s => 
                           key_valid, data_ready_s => key_ready, data_p(31) => 
                           sdi_data(31), data_p(30) => sdi_data(30), data_p(29)
                           => sdi_data(29), data_p(28) => sdi_data(28), 
                           data_p(27) => sdi_data(27), data_p(26) => 
                           sdi_data(26), data_p(25) => sdi_data(25), data_p(24)
                           => sdi_data(24), data_p(23) => sdi_data(23), 
                           data_p(22) => sdi_data(22), data_p(21) => 
                           sdi_data(21), data_p(20) => sdi_data(20), data_p(19)
                           => sdi_data(19), data_p(18) => sdi_data(18), 
                           data_p(17) => sdi_data(17), data_p(16) => 
                           sdi_data(16), data_p(15) => sdi_data(15), data_p(14)
                           => sdi_data(14), data_p(13) => sdi_data(13), 
                           data_p(12) => sdi_data(12), data_p(11) => 
                           sdi_data(11), data_p(10) => sdi_data(10), data_p(9) 
                           => sdi_data(9), data_p(8) => sdi_data(8), data_p(7) 
                           => sdi_data(7), data_p(6) => sdi_data(6), data_p(5) 
                           => sdi_data(5), data_p(4) => sdi_data(4), data_p(3) 
                           => sdi_data(3), data_p(2) => sdi_data(2), data_p(1) 
                           => sdi_data(1), data_p(0) => sdi_data(0), 
                           data_valid_p => key_valid_p, data_ready_p => 
                           key_ready_p);
   bdiPISO : DATA_PISO_1 port map( clk => clk, rst => rst, data_size_p(2) => 
                           bdi_size_p_2_port, data_size_p(1) => 
                           bdi_size_p_1_port, data_size_p(0) => 
                           bdi_size_p_0_port, data_size_s(2) => bdi_size(2), 
                           data_size_s(1) => bdi_size(1), data_size_s(0) => 
                           bdi_size(0), data_s(31) => bdi(31), data_s(30) => 
                           bdi(30), data_s(29) => bdi(29), data_s(28) => 
                           bdi(28), data_s(27) => bdi(27), data_s(26) => 
                           bdi(26), data_s(25) => bdi(25), data_s(24) => 
                           bdi(24), data_s(23) => bdi(23), data_s(22) => 
                           bdi(22), data_s(21) => bdi(21), data_s(20) => 
                           bdi(20), data_s(19) => bdi(19), data_s(18) => 
                           bdi(18), data_s(17) => bdi(17), data_s(16) => 
                           bdi(16), data_s(15) => bdi(15), data_s(14) => 
                           bdi(14), data_s(13) => bdi(13), data_s(12) => 
                           bdi(12), data_s(11) => bdi(11), data_s(10) => 
                           bdi(10), data_s(9) => bdi(9), data_s(8) => bdi(8), 
                           data_s(7) => bdi(7), data_s(6) => bdi(6), data_s(5) 
                           => bdi(5), data_s(4) => bdi(4), data_s(3) => bdi(3),
                           data_s(2) => bdi(2), data_s(1) => bdi(1), data_s(0) 
                           => bdi(0), data_valid_s => bdi_valid, data_ready_s 
                           => bdi_ready, data_p(31) => pdi_data(31), data_p(30)
                           => pdi_data(30), data_p(29) => pdi_data(29), 
                           data_p(28) => pdi_data(28), data_p(27) => 
                           pdi_data(27), data_p(26) => pdi_data(26), data_p(25)
                           => pdi_data(25), data_p(24) => pdi_data(24), 
                           data_p(23) => pdi_data(23), data_p(22) => 
                           pdi_data(22), data_p(21) => pdi_data(21), data_p(20)
                           => pdi_data(20), data_p(19) => pdi_data(19), 
                           data_p(18) => pdi_data(18), data_p(17) => 
                           pdi_data(17), data_p(16) => pdi_data(16), data_p(15)
                           => pdi_data(15), data_p(14) => pdi_data(14), 
                           data_p(13) => pdi_data(13), data_p(12) => 
                           pdi_data(12), data_p(11) => pdi_data(11), data_p(10)
                           => pdi_data(10), data_p(9) => pdi_data(9), data_p(8)
                           => pdi_data(8), data_p(7) => pdi_data(7), data_p(6) 
                           => pdi_data(6), data_p(5) => pdi_data(5), data_p(4) 
                           => pdi_data(4), data_p(3) => pdi_data(3), data_p(2) 
                           => pdi_data(2), data_p(1) => pdi_data(1), data_p(0) 
                           => pdi_data(0), data_valid_p => bdi_valid_p, 
                           data_ready_p => bdi_ready_p, valid_bytes_p(3) => 
                           bdi_valid_bytes_p_3_port, valid_bytes_p(2) => n11, 
                           valid_bytes_p(1) => bdi_valid_bytes_p_1_port, 
                           valid_bytes_p(0) => bdi_valid_bytes_p_0_port, 
                           valid_bytes_s(3) => bdi_valid_bytes(3), 
                           valid_bytes_s(2) => bdi_valid_bytes(2), 
                           valid_bytes_s(1) => bdi_valid_bytes(1), 
                           valid_bytes_s(0) => bdi_valid_bytes(0), pad_loc_p(3)
                           => bdi_pad_loc_p_3_port, pad_loc_p(2) => n14, 
                           pad_loc_p(1) => bdi_pad_loc_p_1_port, pad_loc_p(0) 
                           => bdi_pad_loc_p_0_port, pad_loc_s(3) => 
                           bdi_pad_loc(3), pad_loc_s(2) => bdi_pad_loc(2), 
                           pad_loc_s(1) => bdi_pad_loc(1), pad_loc_s(0) => 
                           bdi_pad_loc(0), eoi_p => bdi_eoi_internal, eoi_s => 
                           bdi_eoi, eot_p => bdi_eot_internal, eot_s => bdi_eot
                           );
   U3 : NAND2X0 port map( IN1 => n52, IN2 => n70, QN => n116);
   U4 : NAND2X0 port map( IN1 => n122, IN2 => n124, QN => n56);
   U5 : NAND2X0 port map( IN1 => n124, IN2 => n103, QN => n53);
   U6 : NOR2X0 port map( IN1 => n27, IN2 => pr_state_2_port, QN => n124);
   U7 : NOR2X0 port map( IN1 => n28, IN2 => pr_state_0_port, QN => n103);
   U8 : NOR2X0 port map( IN1 => n29, IN2 => pr_state_1_port, QN => n114);
   U9 : NOR2X0 port map( IN1 => n28, IN2 => n29, QN => n57);
   U10 : INVX0 port map( INP => n52, ZN => n18);
   U11 : INVX0 port map( INP => n77, ZN => bdi_type_1_port);
   U12 : INVX0 port map( INP => bdi_ready_p, ZN => n7);
   U13 : NOR2X0 port map( IN1 => n19, IN2 => bdi_type_3_port, QN => n52);
   U14 : INVX0 port map( INP => n70, ZN => n21);
   U15 : NOR2X0 port map( IN1 => n22, IN2 => n79, QN => n70);
   U16 : INVX0 port map( INP => n54, ZN => n22);
   U17 : NAND2X1 port map( IN1 => n73, IN2 => n74, QN => bdi_type_3_port);
   U18 : INVX0 port map( INP => n47, ZN => n16);
   U19 : INVX0 port map( INP => n56, ZN => n25);
   U20 : INVX0 port map( INP => n37, ZN => n31);
   U21 : NOR2X0 port map( IN1 => n55, IN2 => n56, QN => n50);
   U22 : INVX0 port map( INP => n38, ZN => n23);
   U23 : INVX0 port map( INP => n72, ZN => n19);
   U24 : INVX0 port map( INP => n76, ZN => n11);
   U25 : INVX0 port map( INP => N64, ZN => n10);
   U26 : NAND2X1 port map( IN1 => n123, IN2 => n114, QN => n73);
   U27 : NAND2X1 port map( IN1 => n124, IN2 => n114, QN => n54);
   U28 : NOR2X0 port map( IN1 => n15, IN2 => n10, QN => bdi_size_p_1_port);
   U29 : NOR2X0 port map( IN1 => n13, IN2 => n10, QN => bdi_size_p_0_port);
   U30 : NAND2X1 port map( IN1 => n124, IN2 => n57, QN => n74);
   U31 : NAND2X0 port map( IN1 => n123, IN2 => n57, QN => n72);
   U32 : INVX0 port map( INP => n104, ZN => n9);
   U33 : INVX0 port map( INP => n87, ZN => n8);
   U34 : NOR2X0 port map( IN1 => n133, IN2 => n65, QN => n90);
   U35 : NOR4X0 port map( IN1 => n50, IN2 => n51, IN3 => n133, IN4 => n18, QN 
                           => n49);
   U36 : NAND2X0 port map( IN1 => n53, IN2 => n54, QN => n51);
   U37 : NOR2X0 port map( IN1 => n133, IN2 => n17, QN => n55);
   U38 : AND2X1 port map( IN1 => n122, IN2 => n110, Q => n41);
   U39 : INVX0 port map( INP => n44, ZN => n26);
   U40 : NAND2X0 port map( IN1 => n123, IN2 => n103, QN => n65);
   U41 : NAND2X0 port map( IN1 => n102, IN2 => n122, QN => n64_port);
   U42 : NAND2X0 port map( IN1 => n122, IN2 => n123, QN => n66);
   U43 : INVX0 port map( INP => n115, ZN => n32);
   U44 : NAND2X1 port map( IN1 => n75, IN2 => n76, QN => 
                           bdi_valid_bytes_p_3_port);
   U45 : NOR2X0 port map( IN1 => bdi_pad_loc_p_1_port, IN2 => 
                           bdi_valid_bytes_p_1_port, QN => n76);
   U46 : INVX0 port map( INP => n60, ZN => n34);
   U47 : NOR4X0 port map( IN1 => bdi_pad_loc_p_1_port, IN2 => n14, IN3 => 
                           bdi_pad_loc_p_3_port, IN4 => bdi_pad_loc_p_0_port, 
                           QN => bdi_valid_bytes_p_0_port);
   U48 : INVX0 port map( INP => n75, ZN => n14);
   U49 : NOR2X0 port map( IN1 => pr_state_3_port, IN2 => pr_state_2_port, QN =>
                           n110);
   U50 : INVX0 port map( INP => dout_SegLenCnt_1_port, ZN => n15);
   U51 : INVX0 port map( INP => dout_SegLenCnt_0_port, ZN => n13);
   U52 : NOR2X0 port map( IN1 => rst, IN2 => n94, QN => N208);
   U53 : NOR2X0 port map( IN1 => rst, IN2 => n98, QN => N207);
   U54 : NOR4X0 port map( IN1 => n99, IN2 => n100, IN3 => n89, IN4 => n97, QN 
                           => n98);
   U55 : NAND2X1 port map( IN1 => n32, IN2 => pdi_valid, QN => n101);
   U56 : INVX0 port map( INP => n65, ZN => n30);
   U57 : NAND2X0 port map( IN1 => n9, IN2 => eot_flag, QN => n87);
   U58 : NAND2X1 port map( IN1 => n109, IN2 => pdi_valid, QN => n108);
   U59 : NOR2X0 port map( IN1 => pr_state_1_port, IN2 => pr_state_0_port, QN =>
                           n122);
   U60 : INVX0 port map( INP => cmd_ready, ZN => n17);
   U61 : NAND3X0 port map( IN1 => sdi_valid, IN2 => key_ready_p, IN3 => N64, QN
                           => n111);
   U62 : NAND3X0 port map( IN1 => n110, IN2 => n111, IN3 => pr_state_1_port, QN
                           => n106);
   U63 : INVX0 port map( INP => n58, ZN => n20);
   U64 : NOR2X0 port map( IN1 => n133, IN2 => n59, QN => n61);
   U65 : NAND2X0 port map( IN1 => n109, IN2 => eot_flag, QN => n115);
   U66 : INVX0 port map( INP => rst, ZN => n33);
   U67 : INVX0 port map( INP => pdi_valid, ZN => n133);
   U68 : INVX0 port map( INP => pdi_data(30), ZN => n36);
   U69 : NOR4X0 port map( IN1 => n125, IN2 => n126, IN3 => n127, IN4 => n128, 
                           QN => n109);
   U70 : NOR4X0 port map( IN1 => n35, IN2 => pdi_data(28), IN3 => pdi_data(29),
                           IN4 => pdi_data(30), QN => n46);
   U71 : NOR4X0 port map( IN1 => dout_SegLenCnt_2_port, IN2 => 
                           dout_SegLenCnt_15_port, IN3 => 
                           dout_SegLenCnt_14_port, IN4 => 
                           dout_SegLenCnt_13_port, QN => n82);
   U72 : NOR4X0 port map( IN1 => dout_SegLenCnt_9_port, IN2 => 
                           dout_SegLenCnt_8_port, IN3 => dout_SegLenCnt_7_port,
                           IN4 => dout_SegLenCnt_6_port, QN => n84);
   U73 : INVX0 port map( INP => pdi_data(31), ZN => n35);
   U74 : INVX0 port map( INP => sdi_valid, ZN => n134);
   U75 : NOR2X0 port map( IN1 => n79, IN2 => n69, QN => n77);
   U76 : AND2X2 port map( IN1 => sdi_valid, IN2 => key_update_port, Q => 
                           key_valid_p);
   U77 : NAND2X0 port map( IN1 => n22, IN2 => decrypt_port, QN => n78);
   U78 : NAND2X0 port map( IN1 => n103, IN2 => n110, QN => n1);
   U113 : NAND2X0 port map( IN1 => n114, IN2 => n110, QN => n38);
   U149 : NAND2X0 port map( IN1 => n103, IN2 => n110, QN => n37);
   U153 : NAND2X0 port map( IN1 => key_ready_p, IN2 => key_update_port, QN => 
                           n39);
   U160 : OA21X1 port map( IN1 => dout_SegLenCnt_0_port, IN2 => 
                           dout_SegLenCnt_1_port, IN3 => dout_SegLenCnt_2_port,
                           Q => n2);
   U171 : NOR3X0 port map( IN1 => n2, IN2 => dout_SegLenCnt_11_port, IN3 => 
                           dout_SegLenCnt_10_port, QN => n6);
   U172 : NOR4X0 port map( IN1 => dout_SegLenCnt_15_port, IN2 => 
                           dout_SegLenCnt_14_port, IN3 => 
                           dout_SegLenCnt_13_port, IN4 => 
                           dout_SegLenCnt_12_port, QN => n5);
   U173 : NOR3X0 port map( IN1 => dout_SegLenCnt_3_port, IN2 => 
                           dout_SegLenCnt_5_port, IN3 => dout_SegLenCnt_4_port,
                           QN => n4);
   U174 : NOR4X0 port map( IN1 => dout_SegLenCnt_9_port, IN2 => 
                           dout_SegLenCnt_8_port, IN3 => dout_SegLenCnt_7_port,
                           IN4 => dout_SegLenCnt_6_port, QN => n3);
   U175 : AND4X1 port map( IN1 => n6, IN2 => n5, IN3 => n4, IN4 => n3, Q => N64
                           );

end SYN_PreProcessor;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_LWC_1.all;

entity LWC_1 is

   port( clk, rst : in std_logic;  pdi_data : in std_logic_vector (31 downto 0)
         ;  pdi_valid : in std_logic;  pdi_ready : out std_logic;  sdi_data : 
         in std_logic_vector (31 downto 0);  sdi_valid : in std_logic;  
         sdi_ready : out std_logic;  do_data : out std_logic_vector (31 downto 
         0);  do_ready : in std_logic;  do_valid, do_last : out std_logic);

end LWC_1;

architecture SYN_structure of LWC_1 is

   component fwft_fifo_G_W32_G_LOG2DEPTH2
      port( clk, rst : in std_logic;  din : in std_logic_vector (31 downto 0); 
            din_valid : in std_logic;  din_ready : out std_logic;  dout : out 
            std_logic_vector (31 downto 0);  dout_valid : out std_logic;  
            dout_ready : in std_logic);
   end component;
   
   component PostProcessor_1
      port( clk, rst : in std_logic;  bdo : in std_logic_vector (31 downto 0); 
            bdo_valid : in std_logic;  bdo_ready : out std_logic;  end_of_block
            : in std_logic;  bdo_type, bdo_valid_bytes : in std_logic_vector (3
            downto 0);  msg_auth : in std_logic;  msg_auth_ready : out 
            std_logic;  msg_auth_valid : in std_logic;  cmd : in 
            std_logic_vector (31 downto 0);  cmd_valid : in std_logic;  
            cmd_ready : out std_logic;  do_data : out std_logic_vector (31 
            downto 0);  do_valid, do_last : out std_logic;  do_ready : in 
            std_logic);
   end component;
   
   component CryptoCore_1
      port( clk, rst : in std_logic;  key : in std_logic_vector (31 downto 0); 
            key_valid : in std_logic;  key_ready : out std_logic;  bdi : in 
            std_logic_vector (31 downto 0);  bdi_valid : in std_logic;  
            bdi_ready : out std_logic;  bdi_pad_loc, bdi_valid_bytes : in 
            std_logic_vector (3 downto 0);  bdi_size : in std_logic_vector (2 
            downto 0);  bdi_eot, bdi_eoi : in std_logic;  bdi_type : in 
            std_logic_vector (3 downto 0);  decrypt_in, key_update, hash_in : 
            in std_logic;  bdo : out std_logic_vector (31 downto 0);  bdo_valid
            : out std_logic;  bdo_ready : in std_logic;  bdo_type, 
            bdo_valid_bytes : out std_logic_vector (3 downto 0);  end_of_block,
            msg_auth_valid : out std_logic;  msg_auth_ready : in std_logic;  
            msg_auth : out std_logic);
   end component;
   
   component PreProcessor_1
      port( clk, rst : in std_logic;  pdi_data : in std_logic_vector (31 downto
            0);  pdi_valid : in std_logic;  pdi_ready : out std_logic;  
            sdi_data : in std_logic_vector (31 downto 0);  sdi_valid : in 
            std_logic;  sdi_ready : out std_logic;  key : out std_logic_vector 
            (31 downto 0);  key_valid : out std_logic;  key_ready : in 
            std_logic;  bdi : out std_logic_vector (31 downto 0);  bdi_valid : 
            out std_logic;  bdi_ready : in std_logic;  bdi_pad_loc, 
            bdi_valid_bytes : out std_logic_vector (3 downto 0);  bdi_size : 
            out std_logic_vector (2 downto 0);  bdi_eot, bdi_eoi : out 
            std_logic;  bdi_type : out std_logic_vector (3 downto 0);  decrypt,
            hash, key_update : out std_logic;  cmd : out std_logic_vector (31 
            downto 0);  cmd_valid : out std_logic;  cmd_ready : in std_logic);
   end component;
   
   signal key_cipher_in_31_port, key_cipher_in_30_port, key_cipher_in_29_port, 
      key_cipher_in_28_port, key_cipher_in_27_port, key_cipher_in_26_port, 
      key_cipher_in_25_port, key_cipher_in_24_port, key_cipher_in_23_port, 
      key_cipher_in_22_port, key_cipher_in_21_port, key_cipher_in_20_port, 
      key_cipher_in_19_port, key_cipher_in_18_port, key_cipher_in_17_port, 
      key_cipher_in_16_port, key_cipher_in_15_port, key_cipher_in_14_port, 
      key_cipher_in_13_port, key_cipher_in_12_port, key_cipher_in_11_port, 
      key_cipher_in_10_port, key_cipher_in_9_port, key_cipher_in_8_port, 
      key_cipher_in_7_port, key_cipher_in_6_port, key_cipher_in_5_port, 
      key_cipher_in_4_port, key_cipher_in_3_port, key_cipher_in_2_port, 
      key_cipher_in_1_port, key_cipher_in_0_port, key_valid_cipher_in, 
      key_ready_cipher_in, bdi_cipher_in_31_port, bdi_cipher_in_30_port, 
      bdi_cipher_in_29_port, bdi_cipher_in_28_port, bdi_cipher_in_27_port, 
      bdi_cipher_in_26_port, bdi_cipher_in_25_port, bdi_cipher_in_24_port, 
      bdi_cipher_in_23_port, bdi_cipher_in_22_port, bdi_cipher_in_21_port, 
      bdi_cipher_in_20_port, bdi_cipher_in_19_port, bdi_cipher_in_18_port, 
      bdi_cipher_in_17_port, bdi_cipher_in_16_port, bdi_cipher_in_15_port, 
      bdi_cipher_in_14_port, bdi_cipher_in_13_port, bdi_cipher_in_12_port, 
      bdi_cipher_in_11_port, bdi_cipher_in_10_port, bdi_cipher_in_9_port, 
      bdi_cipher_in_8_port, bdi_cipher_in_7_port, bdi_cipher_in_6_port, 
      bdi_cipher_in_5_port, bdi_cipher_in_4_port, bdi_cipher_in_3_port, 
      bdi_cipher_in_2_port, bdi_cipher_in_1_port, bdi_cipher_in_0_port, 
      bdi_valid_cipher_in, bdi_ready_cipher_in, bdi_pad_loc_cipher_in_3_port, 
      bdi_pad_loc_cipher_in_2_port, bdi_pad_loc_cipher_in_1_port, 
      bdi_pad_loc_cipher_in_0_port, bdi_valid_bytes_cipher_in_3_port, 
      bdi_valid_bytes_cipher_in_2_port, bdi_valid_bytes_cipher_in_1_port, 
      bdi_valid_bytes_cipher_in_0_port, bdi_size_cipher_in_2_port, 
      bdi_size_cipher_in_1_port, bdi_size_cipher_in_0_port, bdi_eot_cipher_in, 
      bdi_eoi_cipher_in, bdi_type_cipher_in_3_port, bdi_type_cipher_in_2_port, 
      bdi_type_cipher_in_1_port, bdi_type_cipher_in_0_port, decrypt_cipher_in, 
      hash_cipher_in, key_update_cipher_in, cmd_FIFO_in_31_port, 
      cmd_FIFO_in_30_port, cmd_FIFO_in_29_port, cmd_FIFO_in_28_port, 
      cmd_FIFO_in_27_port, cmd_FIFO_in_26_port, cmd_FIFO_in_25_port, 
      cmd_FIFO_in_24_port, cmd_FIFO_in_23_port, cmd_FIFO_in_22_port, 
      cmd_FIFO_in_21_port, cmd_FIFO_in_20_port, cmd_FIFO_in_19_port, 
      cmd_FIFO_in_18_port, cmd_FIFO_in_17_port, cmd_FIFO_in_16_port, 
      cmd_FIFO_in_15_port, cmd_FIFO_in_14_port, cmd_FIFO_in_13_port, 
      cmd_FIFO_in_12_port, cmd_FIFO_in_11_port, cmd_FIFO_in_10_port, 
      cmd_FIFO_in_9_port, cmd_FIFO_in_8_port, cmd_FIFO_in_7_port, 
      cmd_FIFO_in_6_port, cmd_FIFO_in_5_port, cmd_FIFO_in_4_port, 
      cmd_FIFO_in_3_port, cmd_FIFO_in_2_port, cmd_FIFO_in_1_port, 
      cmd_FIFO_in_0_port, cmd_valid_FIFO_in, cmd_ready_FIFO_in, 
      bdo_cipher_out_31_port, bdo_cipher_out_30_port, bdo_cipher_out_29_port, 
      bdo_cipher_out_28_port, bdo_cipher_out_27_port, bdo_cipher_out_26_port, 
      bdo_cipher_out_25_port, bdo_cipher_out_24_port, bdo_cipher_out_23_port, 
      bdo_cipher_out_22_port, bdo_cipher_out_21_port, bdo_cipher_out_20_port, 
      bdo_cipher_out_19_port, bdo_cipher_out_18_port, bdo_cipher_out_17_port, 
      bdo_cipher_out_16_port, bdo_cipher_out_15_port, bdo_cipher_out_14_port, 
      bdo_cipher_out_13_port, bdo_cipher_out_12_port, bdo_cipher_out_11_port, 
      bdo_cipher_out_10_port, bdo_cipher_out_9_port, bdo_cipher_out_8_port, 
      bdo_cipher_out_7_port, bdo_cipher_out_6_port, bdo_cipher_out_5_port, 
      bdo_cipher_out_4_port, bdo_cipher_out_3_port, bdo_cipher_out_2_port, 
      bdo_cipher_out_1_port, bdo_cipher_out_0_port, bdo_valid_cipher_out, 
      bdo_ready_cipher_out, bdo_type_cipher_out_3_port, 
      bdo_type_cipher_out_2_port, bdo_type_cipher_out_1_port, 
      bdo_type_cipher_out_0_port, bdo_valid_bytes_cipher_out_3_port, 
      bdo_valid_bytes_cipher_out_2_port, bdo_valid_bytes_cipher_out_1_port, 
      bdo_valid_bytes_cipher_out_0_port, end_of_block_cipher_out, 
      msg_auth_valid, msg_auth_ready, msg_auth, cmd_FIFO_out_31_port, 
      cmd_FIFO_out_30_port, cmd_FIFO_out_29_port, cmd_FIFO_out_28_port, 
      cmd_FIFO_out_27_port, cmd_FIFO_out_26_port, cmd_FIFO_out_25_port, 
      cmd_FIFO_out_24_port, cmd_FIFO_out_23_port, cmd_FIFO_out_22_port, 
      cmd_FIFO_out_21_port, cmd_FIFO_out_20_port, cmd_FIFO_out_19_port, 
      cmd_FIFO_out_18_port, cmd_FIFO_out_17_port, cmd_FIFO_out_16_port, 
      cmd_FIFO_out_15_port, cmd_FIFO_out_14_port, cmd_FIFO_out_13_port, 
      cmd_FIFO_out_12_port, cmd_FIFO_out_11_port, cmd_FIFO_out_10_port, 
      cmd_FIFO_out_9_port, cmd_FIFO_out_8_port, cmd_FIFO_out_7_port, 
      cmd_FIFO_out_6_port, cmd_FIFO_out_5_port, cmd_FIFO_out_4_port, 
      cmd_FIFO_out_3_port, cmd_FIFO_out_2_port, cmd_FIFO_out_1_port, 
      cmd_FIFO_out_0_port, cmd_valid_FIFO_out, cmd_ready_FIFO_out, n_3235 : 
      std_logic;

begin
   
   Inst_PreProcessor : PreProcessor_1 port map( clk => clk, rst => rst, 
                           pdi_data(31) => pdi_data(31), pdi_data(30) => 
                           pdi_data(30), pdi_data(29) => pdi_data(29), 
                           pdi_data(28) => pdi_data(28), pdi_data(27) => 
                           pdi_data(27), pdi_data(26) => pdi_data(26), 
                           pdi_data(25) => pdi_data(25), pdi_data(24) => 
                           pdi_data(24), pdi_data(23) => pdi_data(23), 
                           pdi_data(22) => pdi_data(22), pdi_data(21) => 
                           pdi_data(21), pdi_data(20) => pdi_data(20), 
                           pdi_data(19) => pdi_data(19), pdi_data(18) => 
                           pdi_data(18), pdi_data(17) => pdi_data(17), 
                           pdi_data(16) => pdi_data(16), pdi_data(15) => 
                           pdi_data(15), pdi_data(14) => pdi_data(14), 
                           pdi_data(13) => pdi_data(13), pdi_data(12) => 
                           pdi_data(12), pdi_data(11) => pdi_data(11), 
                           pdi_data(10) => pdi_data(10), pdi_data(9) => 
                           pdi_data(9), pdi_data(8) => pdi_data(8), pdi_data(7)
                           => pdi_data(7), pdi_data(6) => pdi_data(6), 
                           pdi_data(5) => pdi_data(5), pdi_data(4) => 
                           pdi_data(4), pdi_data(3) => pdi_data(3), pdi_data(2)
                           => pdi_data(2), pdi_data(1) => pdi_data(1), 
                           pdi_data(0) => pdi_data(0), pdi_valid => pdi_valid, 
                           pdi_ready => pdi_ready, sdi_data(31) => sdi_data(31)
                           , sdi_data(30) => sdi_data(30), sdi_data(29) => 
                           sdi_data(29), sdi_data(28) => sdi_data(28), 
                           sdi_data(27) => sdi_data(27), sdi_data(26) => 
                           sdi_data(26), sdi_data(25) => sdi_data(25), 
                           sdi_data(24) => sdi_data(24), sdi_data(23) => 
                           sdi_data(23), sdi_data(22) => sdi_data(22), 
                           sdi_data(21) => sdi_data(21), sdi_data(20) => 
                           sdi_data(20), sdi_data(19) => sdi_data(19), 
                           sdi_data(18) => sdi_data(18), sdi_data(17) => 
                           sdi_data(17), sdi_data(16) => sdi_data(16), 
                           sdi_data(15) => sdi_data(15), sdi_data(14) => 
                           sdi_data(14), sdi_data(13) => sdi_data(13), 
                           sdi_data(12) => sdi_data(12), sdi_data(11) => 
                           sdi_data(11), sdi_data(10) => sdi_data(10), 
                           sdi_data(9) => sdi_data(9), sdi_data(8) => 
                           sdi_data(8), sdi_data(7) => sdi_data(7), sdi_data(6)
                           => sdi_data(6), sdi_data(5) => sdi_data(5), 
                           sdi_data(4) => sdi_data(4), sdi_data(3) => 
                           sdi_data(3), sdi_data(2) => sdi_data(2), sdi_data(1)
                           => sdi_data(1), sdi_data(0) => sdi_data(0), 
                           sdi_valid => sdi_valid, sdi_ready => sdi_ready, 
                           key(31) => key_cipher_in_31_port, key(30) => 
                           key_cipher_in_30_port, key(29) => 
                           key_cipher_in_29_port, key(28) => 
                           key_cipher_in_28_port, key(27) => 
                           key_cipher_in_27_port, key(26) => 
                           key_cipher_in_26_port, key(25) => 
                           key_cipher_in_25_port, key(24) => 
                           key_cipher_in_24_port, key(23) => 
                           key_cipher_in_23_port, key(22) => 
                           key_cipher_in_22_port, key(21) => 
                           key_cipher_in_21_port, key(20) => 
                           key_cipher_in_20_port, key(19) => 
                           key_cipher_in_19_port, key(18) => 
                           key_cipher_in_18_port, key(17) => 
                           key_cipher_in_17_port, key(16) => 
                           key_cipher_in_16_port, key(15) => 
                           key_cipher_in_15_port, key(14) => 
                           key_cipher_in_14_port, key(13) => 
                           key_cipher_in_13_port, key(12) => 
                           key_cipher_in_12_port, key(11) => 
                           key_cipher_in_11_port, key(10) => 
                           key_cipher_in_10_port, key(9) => 
                           key_cipher_in_9_port, key(8) => key_cipher_in_8_port
                           , key(7) => key_cipher_in_7_port, key(6) => 
                           key_cipher_in_6_port, key(5) => key_cipher_in_5_port
                           , key(4) => key_cipher_in_4_port, key(3) => 
                           key_cipher_in_3_port, key(2) => key_cipher_in_2_port
                           , key(1) => key_cipher_in_1_port, key(0) => 
                           key_cipher_in_0_port, key_valid => 
                           key_valid_cipher_in, key_ready => 
                           key_ready_cipher_in, bdi(31) => 
                           bdi_cipher_in_31_port, bdi(30) => 
                           bdi_cipher_in_30_port, bdi(29) => 
                           bdi_cipher_in_29_port, bdi(28) => 
                           bdi_cipher_in_28_port, bdi(27) => 
                           bdi_cipher_in_27_port, bdi(26) => 
                           bdi_cipher_in_26_port, bdi(25) => 
                           bdi_cipher_in_25_port, bdi(24) => 
                           bdi_cipher_in_24_port, bdi(23) => 
                           bdi_cipher_in_23_port, bdi(22) => 
                           bdi_cipher_in_22_port, bdi(21) => 
                           bdi_cipher_in_21_port, bdi(20) => 
                           bdi_cipher_in_20_port, bdi(19) => 
                           bdi_cipher_in_19_port, bdi(18) => 
                           bdi_cipher_in_18_port, bdi(17) => 
                           bdi_cipher_in_17_port, bdi(16) => 
                           bdi_cipher_in_16_port, bdi(15) => 
                           bdi_cipher_in_15_port, bdi(14) => 
                           bdi_cipher_in_14_port, bdi(13) => 
                           bdi_cipher_in_13_port, bdi(12) => 
                           bdi_cipher_in_12_port, bdi(11) => 
                           bdi_cipher_in_11_port, bdi(10) => 
                           bdi_cipher_in_10_port, bdi(9) => 
                           bdi_cipher_in_9_port, bdi(8) => bdi_cipher_in_8_port
                           , bdi(7) => bdi_cipher_in_7_port, bdi(6) => 
                           bdi_cipher_in_6_port, bdi(5) => bdi_cipher_in_5_port
                           , bdi(4) => bdi_cipher_in_4_port, bdi(3) => 
                           bdi_cipher_in_3_port, bdi(2) => bdi_cipher_in_2_port
                           , bdi(1) => bdi_cipher_in_1_port, bdi(0) => 
                           bdi_cipher_in_0_port, bdi_valid => 
                           bdi_valid_cipher_in, bdi_ready => 
                           bdi_ready_cipher_in, bdi_pad_loc(3) => 
                           bdi_pad_loc_cipher_in_3_port, bdi_pad_loc(2) => 
                           bdi_pad_loc_cipher_in_2_port, bdi_pad_loc(1) => 
                           bdi_pad_loc_cipher_in_1_port, bdi_pad_loc(0) => 
                           bdi_pad_loc_cipher_in_0_port, bdi_valid_bytes(3) => 
                           bdi_valid_bytes_cipher_in_3_port, bdi_valid_bytes(2)
                           => bdi_valid_bytes_cipher_in_2_port, 
                           bdi_valid_bytes(1) => 
                           bdi_valid_bytes_cipher_in_1_port, bdi_valid_bytes(0)
                           => bdi_valid_bytes_cipher_in_0_port, bdi_size(2) => 
                           bdi_size_cipher_in_2_port, bdi_size(1) => 
                           bdi_size_cipher_in_1_port, bdi_size(0) => 
                           bdi_size_cipher_in_0_port, bdi_eot => 
                           bdi_eot_cipher_in, bdi_eoi => bdi_eoi_cipher_in, 
                           bdi_type(3) => bdi_type_cipher_in_3_port, 
                           bdi_type(2) => bdi_type_cipher_in_2_port, 
                           bdi_type(1) => bdi_type_cipher_in_1_port, 
                           bdi_type(0) => bdi_type_cipher_in_0_port, decrypt =>
                           decrypt_cipher_in, hash => hash_cipher_in, 
                           key_update => key_update_cipher_in, cmd(31) => 
                           cmd_FIFO_in_31_port, cmd(30) => cmd_FIFO_in_30_port,
                           cmd(29) => cmd_FIFO_in_29_port, cmd(28) => 
                           cmd_FIFO_in_28_port, cmd(27) => cmd_FIFO_in_27_port,
                           cmd(26) => cmd_FIFO_in_26_port, cmd(25) => 
                           cmd_FIFO_in_25_port, cmd(24) => cmd_FIFO_in_24_port,
                           cmd(23) => cmd_FIFO_in_23_port, cmd(22) => 
                           cmd_FIFO_in_22_port, cmd(21) => cmd_FIFO_in_21_port,
                           cmd(20) => cmd_FIFO_in_20_port, cmd(19) => 
                           cmd_FIFO_in_19_port, cmd(18) => cmd_FIFO_in_18_port,
                           cmd(17) => cmd_FIFO_in_17_port, cmd(16) => 
                           cmd_FIFO_in_16_port, cmd(15) => cmd_FIFO_in_15_port,
                           cmd(14) => cmd_FIFO_in_14_port, cmd(13) => 
                           cmd_FIFO_in_13_port, cmd(12) => cmd_FIFO_in_12_port,
                           cmd(11) => cmd_FIFO_in_11_port, cmd(10) => 
                           cmd_FIFO_in_10_port, cmd(9) => cmd_FIFO_in_9_port, 
                           cmd(8) => cmd_FIFO_in_8_port, cmd(7) => 
                           cmd_FIFO_in_7_port, cmd(6) => cmd_FIFO_in_6_port, 
                           cmd(5) => cmd_FIFO_in_5_port, cmd(4) => 
                           cmd_FIFO_in_4_port, cmd(3) => cmd_FIFO_in_3_port, 
                           cmd(2) => cmd_FIFO_in_2_port, cmd(1) => 
                           cmd_FIFO_in_1_port, cmd(0) => cmd_FIFO_in_0_port, 
                           cmd_valid => cmd_valid_FIFO_in, cmd_ready => 
                           cmd_ready_FIFO_in);
   Inst_Cipher : CryptoCore_1 port map( clk => clk, rst => rst, key(31) => 
                           key_cipher_in_31_port, key(30) => 
                           key_cipher_in_30_port, key(29) => 
                           key_cipher_in_29_port, key(28) => 
                           key_cipher_in_28_port, key(27) => 
                           key_cipher_in_27_port, key(26) => 
                           key_cipher_in_26_port, key(25) => 
                           key_cipher_in_25_port, key(24) => 
                           key_cipher_in_24_port, key(23) => 
                           key_cipher_in_23_port, key(22) => 
                           key_cipher_in_22_port, key(21) => 
                           key_cipher_in_21_port, key(20) => 
                           key_cipher_in_20_port, key(19) => 
                           key_cipher_in_19_port, key(18) => 
                           key_cipher_in_18_port, key(17) => 
                           key_cipher_in_17_port, key(16) => 
                           key_cipher_in_16_port, key(15) => 
                           key_cipher_in_15_port, key(14) => 
                           key_cipher_in_14_port, key(13) => 
                           key_cipher_in_13_port, key(12) => 
                           key_cipher_in_12_port, key(11) => 
                           key_cipher_in_11_port, key(10) => 
                           key_cipher_in_10_port, key(9) => 
                           key_cipher_in_9_port, key(8) => key_cipher_in_8_port
                           , key(7) => key_cipher_in_7_port, key(6) => 
                           key_cipher_in_6_port, key(5) => key_cipher_in_5_port
                           , key(4) => key_cipher_in_4_port, key(3) => 
                           key_cipher_in_3_port, key(2) => key_cipher_in_2_port
                           , key(1) => key_cipher_in_1_port, key(0) => 
                           key_cipher_in_0_port, key_valid => 
                           key_valid_cipher_in, key_ready => 
                           key_ready_cipher_in, bdi(31) => 
                           bdi_cipher_in_31_port, bdi(30) => 
                           bdi_cipher_in_30_port, bdi(29) => 
                           bdi_cipher_in_29_port, bdi(28) => 
                           bdi_cipher_in_28_port, bdi(27) => 
                           bdi_cipher_in_27_port, bdi(26) => 
                           bdi_cipher_in_26_port, bdi(25) => 
                           bdi_cipher_in_25_port, bdi(24) => 
                           bdi_cipher_in_24_port, bdi(23) => 
                           bdi_cipher_in_23_port, bdi(22) => 
                           bdi_cipher_in_22_port, bdi(21) => 
                           bdi_cipher_in_21_port, bdi(20) => 
                           bdi_cipher_in_20_port, bdi(19) => 
                           bdi_cipher_in_19_port, bdi(18) => 
                           bdi_cipher_in_18_port, bdi(17) => 
                           bdi_cipher_in_17_port, bdi(16) => 
                           bdi_cipher_in_16_port, bdi(15) => 
                           bdi_cipher_in_15_port, bdi(14) => 
                           bdi_cipher_in_14_port, bdi(13) => 
                           bdi_cipher_in_13_port, bdi(12) => 
                           bdi_cipher_in_12_port, bdi(11) => 
                           bdi_cipher_in_11_port, bdi(10) => 
                           bdi_cipher_in_10_port, bdi(9) => 
                           bdi_cipher_in_9_port, bdi(8) => bdi_cipher_in_8_port
                           , bdi(7) => bdi_cipher_in_7_port, bdi(6) => 
                           bdi_cipher_in_6_port, bdi(5) => bdi_cipher_in_5_port
                           , bdi(4) => bdi_cipher_in_4_port, bdi(3) => 
                           bdi_cipher_in_3_port, bdi(2) => bdi_cipher_in_2_port
                           , bdi(1) => bdi_cipher_in_1_port, bdi(0) => 
                           bdi_cipher_in_0_port, bdi_valid => 
                           bdi_valid_cipher_in, bdi_ready => 
                           bdi_ready_cipher_in, bdi_pad_loc(3) => 
                           bdi_pad_loc_cipher_in_3_port, bdi_pad_loc(2) => 
                           bdi_pad_loc_cipher_in_2_port, bdi_pad_loc(1) => 
                           bdi_pad_loc_cipher_in_1_port, bdi_pad_loc(0) => 
                           bdi_pad_loc_cipher_in_0_port, bdi_valid_bytes(3) => 
                           bdi_valid_bytes_cipher_in_3_port, bdi_valid_bytes(2)
                           => bdi_valid_bytes_cipher_in_2_port, 
                           bdi_valid_bytes(1) => 
                           bdi_valid_bytes_cipher_in_1_port, bdi_valid_bytes(0)
                           => bdi_valid_bytes_cipher_in_0_port, bdi_size(2) => 
                           bdi_size_cipher_in_2_port, bdi_size(1) => 
                           bdi_size_cipher_in_1_port, bdi_size(0) => 
                           bdi_size_cipher_in_0_port, bdi_eot => 
                           bdi_eot_cipher_in, bdi_eoi => bdi_eoi_cipher_in, 
                           bdi_type(3) => bdi_type_cipher_in_3_port, 
                           bdi_type(2) => bdi_type_cipher_in_2_port, 
                           bdi_type(1) => bdi_type_cipher_in_1_port, 
                           bdi_type(0) => bdi_type_cipher_in_0_port, decrypt_in
                           => decrypt_cipher_in, key_update => 
                           key_update_cipher_in, hash_in => hash_cipher_in, 
                           bdo(31) => bdo_cipher_out_31_port, bdo(30) => 
                           bdo_cipher_out_30_port, bdo(29) => 
                           bdo_cipher_out_29_port, bdo(28) => 
                           bdo_cipher_out_28_port, bdo(27) => 
                           bdo_cipher_out_27_port, bdo(26) => 
                           bdo_cipher_out_26_port, bdo(25) => 
                           bdo_cipher_out_25_port, bdo(24) => 
                           bdo_cipher_out_24_port, bdo(23) => 
                           bdo_cipher_out_23_port, bdo(22) => 
                           bdo_cipher_out_22_port, bdo(21) => 
                           bdo_cipher_out_21_port, bdo(20) => 
                           bdo_cipher_out_20_port, bdo(19) => 
                           bdo_cipher_out_19_port, bdo(18) => 
                           bdo_cipher_out_18_port, bdo(17) => 
                           bdo_cipher_out_17_port, bdo(16) => 
                           bdo_cipher_out_16_port, bdo(15) => 
                           bdo_cipher_out_15_port, bdo(14) => 
                           bdo_cipher_out_14_port, bdo(13) => 
                           bdo_cipher_out_13_port, bdo(12) => 
                           bdo_cipher_out_12_port, bdo(11) => 
                           bdo_cipher_out_11_port, bdo(10) => 
                           bdo_cipher_out_10_port, bdo(9) => 
                           bdo_cipher_out_9_port, bdo(8) => 
                           bdo_cipher_out_8_port, bdo(7) => 
                           bdo_cipher_out_7_port, bdo(6) => 
                           bdo_cipher_out_6_port, bdo(5) => 
                           bdo_cipher_out_5_port, bdo(4) => 
                           bdo_cipher_out_4_port, bdo(3) => 
                           bdo_cipher_out_3_port, bdo(2) => 
                           bdo_cipher_out_2_port, bdo(1) => 
                           bdo_cipher_out_1_port, bdo(0) => 
                           bdo_cipher_out_0_port, bdo_valid => 
                           bdo_valid_cipher_out, bdo_ready => 
                           bdo_ready_cipher_out, bdo_type(3) => 
                           bdo_type_cipher_out_3_port, bdo_type(2) => 
                           bdo_type_cipher_out_2_port, bdo_type(1) => n_3235, 
                           bdo_type(0) => bdo_type_cipher_out_0_port, 
                           bdo_valid_bytes(3) => 
                           bdo_valid_bytes_cipher_out_3_port, 
                           bdo_valid_bytes(2) => 
                           bdo_valid_bytes_cipher_out_2_port, 
                           bdo_valid_bytes(1) => 
                           bdo_valid_bytes_cipher_out_1_port, 
                           bdo_valid_bytes(0) => 
                           bdo_valid_bytes_cipher_out_0_port, end_of_block => 
                           end_of_block_cipher_out, msg_auth_valid => 
                           msg_auth_valid, msg_auth_ready => msg_auth_ready, 
                           msg_auth => msg_auth);
   Inst_PostProcessor : PostProcessor_1 port map( clk => clk, rst => rst, 
                           bdo(31) => bdo_cipher_out_31_port, bdo(30) => 
                           bdo_cipher_out_30_port, bdo(29) => 
                           bdo_cipher_out_29_port, bdo(28) => 
                           bdo_cipher_out_28_port, bdo(27) => 
                           bdo_cipher_out_27_port, bdo(26) => 
                           bdo_cipher_out_26_port, bdo(25) => 
                           bdo_cipher_out_25_port, bdo(24) => 
                           bdo_cipher_out_24_port, bdo(23) => 
                           bdo_cipher_out_23_port, bdo(22) => 
                           bdo_cipher_out_22_port, bdo(21) => 
                           bdo_cipher_out_21_port, bdo(20) => 
                           bdo_cipher_out_20_port, bdo(19) => 
                           bdo_cipher_out_19_port, bdo(18) => 
                           bdo_cipher_out_18_port, bdo(17) => 
                           bdo_cipher_out_17_port, bdo(16) => 
                           bdo_cipher_out_16_port, bdo(15) => 
                           bdo_cipher_out_15_port, bdo(14) => 
                           bdo_cipher_out_14_port, bdo(13) => 
                           bdo_cipher_out_13_port, bdo(12) => 
                           bdo_cipher_out_12_port, bdo(11) => 
                           bdo_cipher_out_11_port, bdo(10) => 
                           bdo_cipher_out_10_port, bdo(9) => 
                           bdo_cipher_out_9_port, bdo(8) => 
                           bdo_cipher_out_8_port, bdo(7) => 
                           bdo_cipher_out_7_port, bdo(6) => 
                           bdo_cipher_out_6_port, bdo(5) => 
                           bdo_cipher_out_5_port, bdo(4) => 
                           bdo_cipher_out_4_port, bdo(3) => 
                           bdo_cipher_out_3_port, bdo(2) => 
                           bdo_cipher_out_2_port, bdo(1) => 
                           bdo_cipher_out_1_port, bdo(0) => 
                           bdo_cipher_out_0_port, bdo_valid => 
                           bdo_valid_cipher_out, bdo_ready => 
                           bdo_ready_cipher_out, end_of_block => 
                           end_of_block_cipher_out, bdo_type(3) => 
                           bdo_type_cipher_out_3_port, bdo_type(2) => 
                           bdo_type_cipher_out_2_port, bdo_type(1) => 
                           bdo_type_cipher_out_1_port, bdo_type(0) => 
                           bdo_type_cipher_out_0_port, bdo_valid_bytes(3) => 
                           bdo_valid_bytes_cipher_out_3_port, 
                           bdo_valid_bytes(2) => 
                           bdo_valid_bytes_cipher_out_2_port, 
                           bdo_valid_bytes(1) => 
                           bdo_valid_bytes_cipher_out_1_port, 
                           bdo_valid_bytes(0) => 
                           bdo_valid_bytes_cipher_out_0_port, msg_auth => 
                           msg_auth, msg_auth_ready => msg_auth_ready, 
                           msg_auth_valid => msg_auth_valid, cmd(31) => 
                           cmd_FIFO_out_31_port, cmd(30) => 
                           cmd_FIFO_out_30_port, cmd(29) => 
                           cmd_FIFO_out_29_port, cmd(28) => 
                           cmd_FIFO_out_28_port, cmd(27) => 
                           cmd_FIFO_out_27_port, cmd(26) => 
                           cmd_FIFO_out_26_port, cmd(25) => 
                           cmd_FIFO_out_25_port, cmd(24) => 
                           cmd_FIFO_out_24_port, cmd(23) => 
                           cmd_FIFO_out_23_port, cmd(22) => 
                           cmd_FIFO_out_22_port, cmd(21) => 
                           cmd_FIFO_out_21_port, cmd(20) => 
                           cmd_FIFO_out_20_port, cmd(19) => 
                           cmd_FIFO_out_19_port, cmd(18) => 
                           cmd_FIFO_out_18_port, cmd(17) => 
                           cmd_FIFO_out_17_port, cmd(16) => 
                           cmd_FIFO_out_16_port, cmd(15) => 
                           cmd_FIFO_out_15_port, cmd(14) => 
                           cmd_FIFO_out_14_port, cmd(13) => 
                           cmd_FIFO_out_13_port, cmd(12) => 
                           cmd_FIFO_out_12_port, cmd(11) => 
                           cmd_FIFO_out_11_port, cmd(10) => 
                           cmd_FIFO_out_10_port, cmd(9) => cmd_FIFO_out_9_port,
                           cmd(8) => cmd_FIFO_out_8_port, cmd(7) => 
                           cmd_FIFO_out_7_port, cmd(6) => cmd_FIFO_out_6_port, 
                           cmd(5) => cmd_FIFO_out_5_port, cmd(4) => 
                           cmd_FIFO_out_4_port, cmd(3) => cmd_FIFO_out_3_port, 
                           cmd(2) => cmd_FIFO_out_2_port, cmd(1) => 
                           cmd_FIFO_out_1_port, cmd(0) => cmd_FIFO_out_0_port, 
                           cmd_valid => cmd_valid_FIFO_out, cmd_ready => 
                           cmd_ready_FIFO_out, do_data(31) => do_data(31), 
                           do_data(30) => do_data(30), do_data(29) => 
                           do_data(29), do_data(28) => do_data(28), do_data(27)
                           => do_data(27), do_data(26) => do_data(26), 
                           do_data(25) => do_data(25), do_data(24) => 
                           do_data(24), do_data(23) => do_data(23), do_data(22)
                           => do_data(22), do_data(21) => do_data(21), 
                           do_data(20) => do_data(20), do_data(19) => 
                           do_data(19), do_data(18) => do_data(18), do_data(17)
                           => do_data(17), do_data(16) => do_data(16), 
                           do_data(15) => do_data(15), do_data(14) => 
                           do_data(14), do_data(13) => do_data(13), do_data(12)
                           => do_data(12), do_data(11) => do_data(11), 
                           do_data(10) => do_data(10), do_data(9) => do_data(9)
                           , do_data(8) => do_data(8), do_data(7) => do_data(7)
                           , do_data(6) => do_data(6), do_data(5) => do_data(5)
                           , do_data(4) => do_data(4), do_data(3) => do_data(3)
                           , do_data(2) => do_data(2), do_data(1) => do_data(1)
                           , do_data(0) => do_data(0), do_valid => do_valid, 
                           do_last => do_last, do_ready => do_ready);
   Inst_Header_Fifo : fwft_fifo_G_W32_G_LOG2DEPTH2 port map( clk => clk, rst =>
                           rst, din(31) => cmd_FIFO_in_31_port, din(30) => 
                           cmd_FIFO_in_30_port, din(29) => cmd_FIFO_in_29_port,
                           din(28) => cmd_FIFO_in_28_port, din(27) => 
                           cmd_FIFO_in_27_port, din(26) => cmd_FIFO_in_26_port,
                           din(25) => cmd_FIFO_in_25_port, din(24) => 
                           cmd_FIFO_in_24_port, din(23) => cmd_FIFO_in_23_port,
                           din(22) => cmd_FIFO_in_22_port, din(21) => 
                           cmd_FIFO_in_21_port, din(20) => cmd_FIFO_in_20_port,
                           din(19) => cmd_FIFO_in_19_port, din(18) => 
                           cmd_FIFO_in_18_port, din(17) => cmd_FIFO_in_17_port,
                           din(16) => cmd_FIFO_in_16_port, din(15) => 
                           cmd_FIFO_in_15_port, din(14) => cmd_FIFO_in_14_port,
                           din(13) => cmd_FIFO_in_13_port, din(12) => 
                           cmd_FIFO_in_12_port, din(11) => cmd_FIFO_in_11_port,
                           din(10) => cmd_FIFO_in_10_port, din(9) => 
                           cmd_FIFO_in_9_port, din(8) => cmd_FIFO_in_8_port, 
                           din(7) => cmd_FIFO_in_7_port, din(6) => 
                           cmd_FIFO_in_6_port, din(5) => cmd_FIFO_in_5_port, 
                           din(4) => cmd_FIFO_in_4_port, din(3) => 
                           cmd_FIFO_in_3_port, din(2) => cmd_FIFO_in_2_port, 
                           din(1) => cmd_FIFO_in_1_port, din(0) => 
                           cmd_FIFO_in_0_port, din_valid => cmd_valid_FIFO_in, 
                           din_ready => cmd_ready_FIFO_in, dout(31) => 
                           cmd_FIFO_out_31_port, dout(30) => 
                           cmd_FIFO_out_30_port, dout(29) => 
                           cmd_FIFO_out_29_port, dout(28) => 
                           cmd_FIFO_out_28_port, dout(27) => 
                           cmd_FIFO_out_27_port, dout(26) => 
                           cmd_FIFO_out_26_port, dout(25) => 
                           cmd_FIFO_out_25_port, dout(24) => 
                           cmd_FIFO_out_24_port, dout(23) => 
                           cmd_FIFO_out_23_port, dout(22) => 
                           cmd_FIFO_out_22_port, dout(21) => 
                           cmd_FIFO_out_21_port, dout(20) => 
                           cmd_FIFO_out_20_port, dout(19) => 
                           cmd_FIFO_out_19_port, dout(18) => 
                           cmd_FIFO_out_18_port, dout(17) => 
                           cmd_FIFO_out_17_port, dout(16) => 
                           cmd_FIFO_out_16_port, dout(15) => 
                           cmd_FIFO_out_15_port, dout(14) => 
                           cmd_FIFO_out_14_port, dout(13) => 
                           cmd_FIFO_out_13_port, dout(12) => 
                           cmd_FIFO_out_12_port, dout(11) => 
                           cmd_FIFO_out_11_port, dout(10) => 
                           cmd_FIFO_out_10_port, dout(9) => cmd_FIFO_out_9_port
                           , dout(8) => cmd_FIFO_out_8_port, dout(7) => 
                           cmd_FIFO_out_7_port, dout(6) => cmd_FIFO_out_6_port,
                           dout(5) => cmd_FIFO_out_5_port, dout(4) => 
                           cmd_FIFO_out_4_port, dout(3) => cmd_FIFO_out_3_port,
                           dout(2) => cmd_FIFO_out_2_port, dout(1) => 
                           cmd_FIFO_out_1_port, dout(0) => cmd_FIFO_out_0_port,
                           dout_valid => cmd_valid_FIFO_out, dout_ready => 
                           cmd_ready_FIFO_out);
   bdo_type_cipher_out_1_port <= '0';

end SYN_structure;
