
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_LWC_1 is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_LWC_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_LWC_1.all;

entity xoodoo_round_ADDRESS_LEN384_1 is

   port( INPUT : in std_logic_vector (383 downto 0);  perm_output : out 
         std_logic_vector (383 downto 0);  RNDCTR : in std_logic_vector (3 
         downto 0));

end xoodoo_round_ADDRESS_LEN384_1;

architecture SYN_Behavioral of xoodoo_round_ADDRESS_LEN384_1 is

   component GTECH_XOR2
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component GTECH_AND2
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component GTECH_NOT
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component SELECT_OP
      generic( num_inputs, input_width : integer );
      port( DATA : in std_logic_vector( num_inputs* input_width - 1 downto 0 );
            CONTROL : in std_logic_vector( num_inputs - 1 downto 0 ); Z : out 
            std_logic_vector( input_width - 1 downto 0 ) );
   end component;
   
   component GTECH_BUF
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component GTECH_AND3
      port( A, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component GTECH_AND4
      port( A, B, C, D : in std_logic;  Z : out std_logic);
   end component;
   
   signal N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15,
      N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30
      , N31, X_Logic1_port, X_Logic0_port, N32, N33, N34, N35, N36, N37, N38, 
      N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53
      , N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, 
      N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82
      , N83, N84, N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, 
      N97, N98, N99, N100, N101, N102, N103, N104, N105, N106, N107, N108, N109
      , N110, N111, N112, N113, N114, N115, N116, N117, N118, N119, N120, N121,
      N122, N123, N124, N125, N126, N127, N128, N129, N130, N131, N132, N133, 
      N134, N135, N136, N137, N138, N139, N140, N141, N142, N143, N144, N145, 
      N146, N147, N148, N149, N150, N151, N152, N153, N154, N155, N156, N157, 
      N158, N159, p_plane_127_port, p_plane_126_port, p_plane_125_port, 
      p_plane_124_port, p_plane_123_port, p_plane_122_port, p_plane_121_port, 
      p_plane_120_port, p_plane_119_port, p_plane_118_port, p_plane_117_port, 
      p_plane_116_port, p_plane_115_port, p_plane_114_port, p_plane_113_port, 
      p_plane_112_port, p_plane_111_port, p_plane_110_port, p_plane_109_port, 
      p_plane_108_port, p_plane_107_port, p_plane_106_port, p_plane_105_port, 
      p_plane_104_port, p_plane_103_port, p_plane_102_port, p_plane_101_port, 
      p_plane_100_port, p_plane_99_port, p_plane_98_port, p_plane_97_port, 
      p_plane_96_port, p_plane_95_port, p_plane_94_port, p_plane_93_port, 
      p_plane_92_port, p_plane_91_port, p_plane_90_port, p_plane_89_port, 
      p_plane_88_port, p_plane_87_port, p_plane_86_port, p_plane_85_port, 
      p_plane_84_port, p_plane_83_port, p_plane_82_port, p_plane_81_port, 
      p_plane_80_port, p_plane_79_port, p_plane_78_port, p_plane_77_port, 
      p_plane_76_port, p_plane_75_port, p_plane_74_port, p_plane_73_port, 
      p_plane_72_port, p_plane_71_port, p_plane_70_port, p_plane_69_port, 
      p_plane_68_port, p_plane_67_port, p_plane_66_port, p_plane_65_port, 
      p_plane_64_port, p_plane_63_port, p_plane_62_port, p_plane_61_port, 
      p_plane_60_port, p_plane_59_port, p_plane_58_port, p_plane_57_port, 
      p_plane_56_port, p_plane_55_port, p_plane_54_port, p_plane_53_port, 
      p_plane_52_port, p_plane_51_port, p_plane_50_port, p_plane_49_port, 
      p_plane_48_port, p_plane_47_port, p_plane_46_port, p_plane_45_port, 
      p_plane_44_port, p_plane_43_port, p_plane_42_port, p_plane_41_port, 
      p_plane_40_port, p_plane_39_port, p_plane_38_port, p_plane_37_port, 
      p_plane_36_port, p_plane_35_port, p_plane_34_port, p_plane_33_port, 
      p_plane_32_port, p_plane_31_port, p_plane_30_port, p_plane_29_port, 
      p_plane_28_port, p_plane_27_port, p_plane_26_port, p_plane_25_port, 
      p_plane_24_port, p_plane_23_port, p_plane_22_port, p_plane_21_port, 
      p_plane_20_port, p_plane_19_port, p_plane_18_port, p_plane_17_port, 
      p_plane_16_port, p_plane_15_port, p_plane_14_port, p_plane_13_port, 
      p_plane_12_port, p_plane_11_port, p_plane_10_port, p_plane_9_port, 
      p_plane_8_port, p_plane_7_port, p_plane_6_port, p_plane_5_port, 
      p_plane_4_port, p_plane_3_port, p_plane_2_port, p_plane_1_port, 
      p_plane_0_port, eshift_127_port, eshift_126_port, eshift_125_port, 
      eshift_124_port, eshift_123_port, eshift_122_port, eshift_121_port, 
      eshift_120_port, eshift_119_port, eshift_118_port, eshift_117_port, 
      eshift_116_port, eshift_115_port, eshift_114_port, eshift_113_port, 
      eshift_112_port, eshift_111_port, eshift_110_port, eshift_109_port, 
      eshift_108_port, eshift_107_port, eshift_106_port, eshift_105_port, 
      eshift_104_port, eshift_103_port, eshift_102_port, eshift_101_port, 
      eshift_100_port, eshift_99_port, eshift_98_port, eshift_97_port, 
      eshift_96_port, eshift_95_port, eshift_94_port, eshift_93_port, 
      eshift_92_port, eshift_91_port, eshift_90_port, eshift_89_port, 
      eshift_88_port, eshift_87_port, eshift_86_port, eshift_85_port, 
      eshift_84_port, eshift_83_port, eshift_82_port, eshift_81_port, 
      eshift_80_port, eshift_79_port, eshift_78_port, eshift_77_port, 
      eshift_76_port, eshift_75_port, eshift_74_port, eshift_73_port, 
      eshift_72_port, eshift_71_port, eshift_70_port, eshift_69_port, 
      eshift_68_port, eshift_67_port, eshift_66_port, eshift_65_port, 
      eshift_64_port, eshift_63_port, eshift_62_port, eshift_61_port, 
      eshift_60_port, eshift_59_port, eshift_58_port, eshift_57_port, 
      eshift_56_port, eshift_55_port, eshift_54_port, eshift_53_port, 
      eshift_52_port, eshift_51_port, eshift_50_port, eshift_49_port, 
      eshift_48_port, eshift_47_port, eshift_46_port, eshift_45_port, 
      eshift_44_port, eshift_43_port, eshift_42_port, eshift_41_port, 
      eshift_40_port, eshift_39_port, eshift_38_port, eshift_37_port, 
      eshift_36_port, eshift_35_port, eshift_34_port, eshift_33_port, 
      eshift_32_port, eshift_31_port, eshift_30_port, eshift_29_port, 
      eshift_28_port, eshift_27_port, eshift_26_port, eshift_25_port, 
      eshift_24_port, eshift_23_port, eshift_22_port, eshift_21_port, 
      eshift_20_port, eshift_19_port, eshift_18_port, eshift_17_port, 
      eshift_16_port, eshift_15_port, eshift_14_port, eshift_13_port, 
      eshift_12_port, eshift_11_port, eshift_10_port, eshift_9_port, 
      eshift_8_port, eshift_7_port, eshift_6_port, eshift_5_port, eshift_4_port
      , eshift_3_port, eshift_2_port, eshift_1_port, eshift_0_port, 
      plane2_2_127_port, plane2_2_126_port, plane2_2_125_port, 
      plane2_2_124_port, plane2_2_123_port, plane2_2_122_port, 
      plane2_2_121_port, plane2_2_120_port, plane2_2_119_port, 
      plane2_2_118_port, plane2_2_117_port, plane2_2_116_port, 
      plane2_2_115_port, plane2_2_114_port, plane2_2_113_port, 
      plane2_2_112_port, plane2_2_111_port, plane2_2_110_port, 
      plane2_2_109_port, plane2_2_108_port, plane2_2_107_port, 
      plane2_2_106_port, plane2_2_105_port, plane2_2_104_port, 
      plane2_2_103_port, plane2_2_102_port, plane2_2_101_port, 
      plane2_2_100_port, plane2_2_99_port, plane2_2_98_port, plane2_2_97_port, 
      plane2_2_96_port, plane2_2_95_port, plane2_2_94_port, plane2_2_93_port, 
      plane2_2_92_port, plane2_2_91_port, plane2_2_90_port, plane2_2_89_port, 
      plane2_2_88_port, plane2_2_87_port, plane2_2_86_port, plane2_2_85_port, 
      plane2_2_84_port, plane2_2_83_port, plane2_2_82_port, plane2_2_81_port, 
      plane2_2_80_port, plane2_2_79_port, plane2_2_78_port, plane2_2_77_port, 
      plane2_2_76_port, plane2_2_75_port, plane2_2_74_port, plane2_2_73_port, 
      plane2_2_72_port, plane2_2_71_port, plane2_2_70_port, plane2_2_69_port, 
      plane2_2_68_port, plane2_2_67_port, plane2_2_66_port, plane2_2_65_port, 
      plane2_2_64_port, plane2_2_63_port, plane2_2_62_port, plane2_2_61_port, 
      plane2_2_60_port, plane2_2_59_port, plane2_2_58_port, plane2_2_57_port, 
      plane2_2_56_port, plane2_2_55_port, plane2_2_54_port, plane2_2_53_port, 
      plane2_2_52_port, plane2_2_51_port, plane2_2_50_port, plane2_2_49_port, 
      plane2_2_48_port, plane2_2_47_port, plane2_2_46_port, plane2_2_45_port, 
      plane2_2_44_port, plane2_2_43_port, plane2_2_42_port, plane2_2_41_port, 
      plane2_2_40_port, plane2_2_39_port, plane2_2_38_port, plane2_2_37_port, 
      plane2_2_36_port, plane2_2_35_port, plane2_2_34_port, plane2_2_33_port, 
      plane2_2_32_port, plane2_2_31_port, plane2_2_30_port, plane2_2_29_port, 
      plane2_2_28_port, plane2_2_27_port, plane2_2_26_port, plane2_2_25_port, 
      plane2_2_24_port, plane2_2_23_port, plane2_2_22_port, plane2_2_21_port, 
      plane2_2_20_port, plane2_2_19_port, plane2_2_18_port, plane2_2_17_port, 
      plane2_2_16_port, plane2_2_15_port, plane2_2_14_port, plane2_2_13_port, 
      plane2_2_12_port, plane2_2_11_port, plane2_2_10_port, plane2_2_9_port, 
      plane2_2_8_port, plane2_2_7_port, plane2_2_6_port, plane2_2_5_port, 
      plane2_2_4_port, plane2_2_3_port, plane2_2_2_port, plane2_2_1_port, 
      plane2_2_0_port, plane1_2_127_port, plane1_2_126_port, plane1_2_125_port,
      plane1_2_124_port, plane1_2_123_port, plane1_2_122_port, 
      plane1_2_121_port, plane1_2_120_port, plane1_2_119_port, 
      plane1_2_118_port, plane1_2_117_port, plane1_2_116_port, 
      plane1_2_115_port, plane1_2_114_port, plane1_2_113_port, 
      plane1_2_112_port, plane1_2_111_port, plane1_2_110_port, 
      plane1_2_109_port, plane1_2_108_port, plane1_2_107_port, 
      plane1_2_106_port, plane1_2_105_port, plane1_2_104_port, 
      plane1_2_103_port, plane1_2_102_port, plane1_2_101_port, 
      plane1_2_100_port, plane1_2_99_port, plane1_2_98_port, plane1_2_97_port, 
      plane1_2_96_port, plane1_2_95_port, plane1_2_94_port, plane1_2_93_port, 
      plane1_2_92_port, plane1_2_91_port, plane1_2_90_port, plane1_2_89_port, 
      plane1_2_88_port, plane1_2_87_port, plane1_2_86_port, plane1_2_85_port, 
      plane1_2_84_port, plane1_2_83_port, plane1_2_82_port, plane1_2_81_port, 
      plane1_2_80_port, plane1_2_79_port, plane1_2_78_port, plane1_2_77_port, 
      plane1_2_76_port, plane1_2_75_port, plane1_2_74_port, plane1_2_73_port, 
      plane1_2_72_port, plane1_2_71_port, plane1_2_70_port, plane1_2_69_port, 
      plane1_2_68_port, plane1_2_67_port, plane1_2_66_port, plane1_2_65_port, 
      plane1_2_64_port, plane1_2_63_port, plane1_2_62_port, plane1_2_61_port, 
      plane1_2_60_port, plane1_2_59_port, plane1_2_58_port, plane1_2_57_port, 
      plane1_2_56_port, plane1_2_55_port, plane1_2_54_port, plane1_2_53_port, 
      plane1_2_52_port, plane1_2_51_port, plane1_2_50_port, plane1_2_49_port, 
      plane1_2_48_port, plane1_2_47_port, plane1_2_46_port, plane1_2_45_port, 
      plane1_2_44_port, plane1_2_43_port, plane1_2_42_port, plane1_2_41_port, 
      plane1_2_40_port, plane1_2_39_port, plane1_2_38_port, plane1_2_37_port, 
      plane1_2_36_port, plane1_2_35_port, plane1_2_34_port, plane1_2_33_port, 
      plane1_2_32_port, plane1_2_31_port, plane1_2_30_port, plane1_2_29_port, 
      plane1_2_28_port, plane1_2_27_port, plane1_2_26_port, plane1_2_25_port, 
      plane1_2_24_port, plane1_2_23_port, plane1_2_22_port, plane1_2_21_port, 
      plane1_2_20_port, plane1_2_19_port, plane1_2_18_port, plane1_2_17_port, 
      plane1_2_16_port, plane1_2_15_port, plane1_2_14_port, plane1_2_13_port, 
      plane1_2_12_port, plane1_2_11_port, plane1_2_10_port, plane1_2_9_port, 
      plane1_2_8_port, plane1_2_7_port, plane1_2_6_port, plane1_2_5_port, 
      plane1_2_4_port, plane1_2_3_port, plane1_2_2_port, plane1_2_1_port, 
      plane1_2_0_port, plane0_2_127_port, plane0_2_126_port, plane0_2_125_port,
      plane0_2_124_port, plane0_2_123_port, plane0_2_122_port, 
      plane0_2_121_port, plane0_2_120_port, plane0_2_119_port, 
      plane0_2_118_port, plane0_2_117_port, plane0_2_116_port, 
      plane0_2_115_port, plane0_2_114_port, plane0_2_113_port, 
      plane0_2_112_port, plane0_2_111_port, plane0_2_110_port, 
      plane0_2_109_port, plane0_2_108_port, plane0_2_107_port, 
      plane0_2_106_port, plane0_2_105_port, plane0_2_104_port, 
      plane0_2_103_port, plane0_2_102_port, plane0_2_101_port, 
      plane0_2_100_port, plane0_2_99_port, plane0_2_98_port, plane0_2_97_port, 
      plane0_2_96_port, plane0_2_95_port, plane0_2_94_port, plane0_2_93_port, 
      plane0_2_92_port, plane0_2_91_port, plane0_2_90_port, plane0_2_89_port, 
      plane0_2_88_port, plane0_2_87_port, plane0_2_86_port, plane0_2_85_port, 
      plane0_2_84_port, plane0_2_83_port, plane0_2_82_port, plane0_2_81_port, 
      plane0_2_80_port, plane0_2_79_port, plane0_2_78_port, plane0_2_77_port, 
      plane0_2_76_port, plane0_2_75_port, plane0_2_74_port, plane0_2_73_port, 
      plane0_2_72_port, plane0_2_71_port, plane0_2_70_port, plane0_2_69_port, 
      plane0_2_68_port, plane0_2_67_port, plane0_2_66_port, plane0_2_65_port, 
      plane0_2_64_port, plane0_2_63_port, plane0_2_62_port, plane0_2_61_port, 
      plane0_2_60_port, plane0_2_59_port, plane0_2_58_port, plane0_2_57_port, 
      plane0_2_56_port, plane0_2_55_port, plane0_2_54_port, plane0_2_53_port, 
      plane0_2_52_port, plane0_2_51_port, plane0_2_50_port, plane0_2_49_port, 
      plane0_2_48_port, plane0_2_47_port, plane0_2_46_port, plane0_2_45_port, 
      plane0_2_44_port, plane0_2_43_port, plane0_2_42_port, plane0_2_41_port, 
      plane0_2_40_port, plane0_2_39_port, plane0_2_38_port, plane0_2_37_port, 
      plane0_2_36_port, plane0_2_35_port, plane0_2_34_port, plane0_2_33_port, 
      plane0_2_32_port, plane0_2_31_port, plane0_2_30_port, plane0_2_29_port, 
      plane0_2_28_port, plane0_2_27_port, plane0_2_26_port, plane0_2_25_port, 
      plane0_2_24_port, plane0_2_23_port, plane0_2_22_port, plane0_2_21_port, 
      plane0_2_20_port, plane0_2_19_port, plane0_2_18_port, plane0_2_17_port, 
      plane0_2_16_port, plane0_2_15_port, plane0_2_14_port, plane0_2_13_port, 
      plane0_2_12_port, plane0_2_11_port, plane0_2_10_port, plane0_2_9_port, 
      plane0_2_8_port, plane0_2_7_port, plane0_2_6_port, plane0_2_5_port, 
      plane0_2_4_port, plane0_2_3_port, plane0_2_2_port, plane0_2_1_port, 
      plane0_2_0_port, N160, N161, N162, N163, N164, N165, N166, N167, N168, 
      N169, N170, N171, N172, N173, N174, N175, N176, N177, N178, N179, N180, 
      add_rnd_const_small_11_port, add_rnd_const_small_10_port, 
      add_rnd_const_small_9_port, add_rnd_const_small_8_port, 
      add_rnd_const_small_7_port, add_rnd_const_small_6_port, 
      add_rnd_const_small_5_port, add_rnd_const_small_4_port, 
      add_rnd_const_small_3_port, add_rnd_const_small_2_port, 
      add_rnd_const_small_1_port, add_rnd_const_small_0_port, N181, N182, N183,
      N184, N185, N186, N187, N188, N189, N190, N191, N192, N193, N194, N195, 
      N196, N197, N198, N199, N200, N201, N202, N203, N204, N205, N206, N207, 
      N208, N209, N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, 
      N220, N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231, 
      N232, N233, N234, N235, N236, N237, N238, N239, N240, N241, N242, N243, 
      N244, N245, N246, N247, N248, N249, N250, N251, N252, N253, N254, N255, 
      N256, N257, N258, N259, N260, N261, N262, N263, N264, N265, N266, N267, 
      N268, N269, N270, N271, N272, N273, N274, N275, N276, N277, N278, N279, 
      N280, N281, N282, N283, N284, N285, N286, N287, N288, N289, N290, N291, 
      N292, N293, N294, N295, N296, N297, N298, N299, N300, N301, N302, N303, 
      N304, N305, N306, N307, N308, N309, N310, N311, N312, N313, N314, N315, 
      N316, N317, N318, N319, N320, N321, N322, N323, N324, N325, N326, N327, 
      N328, N329, N330, N331, N332, N333, N334, N335, N336, N337, N338, N339, 
      N340, N341, N342, N343, N344, N345, N346, N347, N348, N349, N350, N351, 
      N352, N353, N354, N355, N356, N357, N358, N359, N360, N361, N362, N363, 
      N364, N365, N366, N367, N368, N369, N370, N371, N372, N373, N374, N375, 
      N376, N377, N378, N379, N380, N381, N382, N383, N384, N385, N386, N387, 
      N388, N389, N390, N391, N392, N393, N394, N395, N396, N397, N398, N399, 
      N400, N401, N402, N403, N404, N405, N406, N407, N408, N409, N410, N411, 
      N412, N413, N414, N415, N416, N417, N418, N419, N420, N421, N422, N423, 
      N424, N425, N426, N427, N428, N429, N430, N431, N432, N433, N434, N435, 
      N436, N437, N438, N439, N440, N441, N442, N443, N444, N445, N446, N447, 
      N448, N449, N450, N451, N452, N453, N454, N455, N456, N457, N458, N459, 
      N460, N461, N462, N463, N464, N465, N466, N467, N468, N469, N470, N471, 
      N472, N473, N474, N475, N476, N477, N478, N479, N480, N481, N482, N483, 
      N484, N485, N486, N487, N488, N489, N490, N491, N492, N493, N494, N495, 
      N496, N497, N498, N499, N500, N501, N502, N503, N504, N505, N506, N507, 
      N508, N509, N510, N511, N512, N513, N514, N515, N516, N517, N518, N519, 
      N520, N521, N522, N523, N524, N525, N526, N527, N528, N529, N530, N531, 
      N532, N533, N534, N535, N536, N537, N538, N539, N540, N541, N542, N543, 
      N544, N545, N546, N547, N548, N549, N550, N551, N552, N553, N554, N555, 
      N556, N557, N558, N559, N560, N561, N562, N563, N564, N565, N566, N567, 
      N568, N569, N570, N571, N572, N573, N574, N575, N576, N577, N578, N579, 
      N580, N581, N582, N583, N584, N585, N586, N587, N588, N589, N590, N591, 
      N592, N593, N594, N595, N596, N597, N598, N599, N600, N601, N602, N603, 
      N604, N605, N606, N607, N608, N609, N610, N611, N612, N613, N614, N615, 
      N616, N617, N618, N619, N620, N621, N622, N623, N624, N625, N626, N627, 
      N628, N629, N630, N631, N632, N633, N634, N635, N636, N637, N638, N639, 
      N640, N641, N642, N643, N644, N645, N646, N647, N648, N649, N650, N651, 
      N652, N653, N654, N655, N656, N657, N658, N659, N660, N661, N662, N663, 
      N664, N665, N666, N667, N668, N669, N670, N671, N672, N673, N674, N675, 
      N676, N677, N678, N679, N680, N681, N682, N683, N684, N685, N686, N687, 
      N688, N689, N690, N691, N692, N693, N694, N695, N696, N697, N698, N699, 
      N700, N701, N702, N703, N704, N705, N706, N707, N708, N709, N710, N711, 
      N712, N713, N714, N715, N716, N717, N718, N719, N720, N721, N722, N723, 
      N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, 
      N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, 
      N748, N749, N750, N751, N752, N753, N754, N755, N756, N757, N758, N759, 
      N760, N761, N762, N763, N764, N765, N766, N767, N768, N769, N770, N771, 
      N772, N773, N774, N775, N776, N777, N778, N779, N780, N781, N782, N783, 
      N784, N785, N786, N787, N788, N789, N790, N791, N792, N793, N794, N795, 
      N796, N797, N798, N799, N800, N801, N802, N803, N804, N805, N806, N807, 
      N808, N809, N810, N811, N812, N813, N814, N815, N816, N817, N818, N819, 
      N820, N821, N822, N823, N824, N825, N826, N827, N828, N829, N830, N831, 
      N832, N833, N834, N835, N836, N837, N838, N839, N840, N841, N842, N843, 
      N844, N845, N846, N847, N848, N849, N850, N851, N852, N853, N854, N855, 
      N856, N857, N858, N859, N860, N861, N862, N863, N864, N865, N866, N867, 
      N868, N869, N870, N871, N872, N873, N874, N875, N876, N877, N878, N879, 
      N880, N881, N882, N883, N884, N885, N886, N887, N888, N889, N890, N891, 
      N892, N893, N894, N895, N896, N897, N898, N899, N900, N901, N902, N903, 
      N904, N905, N906, N907, N908, N909, N910, N911, N912, N913, N914, N915, 
      N916, N917, N918, N919, N920, N921, N922, N923, N924, N925, N926, N927, 
      N928, N929, N930, N931, N932, N933, N934, N935, N936, N937, N938, N939, 
      N940, N941, N942, N943, N944, N945, N946, N947, N948 : std_logic;

begin
   
   C1990 : GTECH_AND4 port map( A => N0, B => N1, C => N2, D => N3, Z => N160);
   I_0 : GTECH_NOT port map( A => RNDCTR(3), Z => N0);
   I_1 : GTECH_NOT port map( A => RNDCTR(2), Z => N1);
   I_2 : GTECH_NOT port map( A => RNDCTR(0), Z => N2);
   I_3 : GTECH_NOT port map( A => RNDCTR(1), Z => N3);
   C1991 : GTECH_AND3 port map( A => RNDCTR(3), B => N4, C => N5, Z => N161);
   I_4 : GTECH_NOT port map( A => RNDCTR(0), Z => N4);
   I_5 : GTECH_NOT port map( A => RNDCTR(1), Z => N5);
   C1992 : GTECH_AND4 port map( A => N6, B => N7, C => RNDCTR(0), D => N8, Z =>
                           N162);
   I_6 : GTECH_NOT port map( A => RNDCTR(3), Z => N6);
   I_7 : GTECH_NOT port map( A => RNDCTR(2), Z => N7);
   I_8 : GTECH_NOT port map( A => RNDCTR(1), Z => N8);
   C1993 : GTECH_AND4 port map( A => N9, B => N10, C => N11, D => RNDCTR(1), Z 
                           => N164);
   I_9 : GTECH_NOT port map( A => RNDCTR(3), Z => N9);
   I_10 : GTECH_NOT port map( A => RNDCTR(2), Z => N10);
   I_11 : GTECH_NOT port map( A => RNDCTR(0), Z => N11);
   C1994 : GTECH_AND4 port map( A => N12, B => N13, C => RNDCTR(0), D => 
                           RNDCTR(1), Z => N166);
   I_12 : GTECH_NOT port map( A => RNDCTR(3), Z => N12);
   I_13 : GTECH_NOT port map( A => RNDCTR(2), Z => N13);
   C1995 : GTECH_AND3 port map( A => RNDCTR(2), B => N14, C => N15, Z => N168);
   I_14 : GTECH_NOT port map( A => RNDCTR(0), Z => N14);
   I_15 : GTECH_NOT port map( A => RNDCTR(1), Z => N15);
   C1996 : GTECH_AND3 port map( A => RNDCTR(2), B => RNDCTR(0), C => N16, Z => 
                           N169);
   I_16 : GTECH_NOT port map( A => RNDCTR(1), Z => N16);
   C1997 : GTECH_AND3 port map( A => RNDCTR(2), B => N17, C => RNDCTR(1), Z => 
                           N170);
   I_17 : GTECH_NOT port map( A => RNDCTR(0), Z => N17);
   C1998 : GTECH_AND3 port map( A => RNDCTR(2), B => RNDCTR(0), C => RNDCTR(1),
                           Z => N171);
   C1999 : GTECH_AND3 port map( A => RNDCTR(3), B => RNDCTR(0), C => N18, Z => 
                           N163);
   I_18 : GTECH_NOT port map( A => RNDCTR(1), Z => N18);
   C2000 : GTECH_AND3 port map( A => RNDCTR(3), B => N19, C => RNDCTR(1), Z => 
                           N165);
   I_19 : GTECH_NOT port map( A => RNDCTR(0), Z => N19);
   C2001 : GTECH_AND3 port map( A => RNDCTR(3), B => RNDCTR(0), C => RNDCTR(1),
                           Z => N167);
   C2006_cell : SELECT_OP
      generic map ( num_inputs => 12, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => X_Logic0_port, 
         -- Connections to port 'DATA3'
         DATA(2) => X_Logic1_port, 
         -- Connections to port 'DATA4'
         DATA(3) => X_Logic0_port, 
         -- Connections to port 'DATA5'
         DATA(4) => X_Logic0_port, 
         -- Connections to port 'DATA6'
         DATA(5) => X_Logic0_port, 
         -- Connections to port 'DATA7'
         DATA(6) => X_Logic0_port, 
         -- Connections to port 'DATA8'
         DATA(7) => X_Logic0_port, 
         -- Connections to port 'DATA9'
         DATA(8) => X_Logic1_port, 
         -- Connections to port 'DATA10'
         DATA(9) => X_Logic0_port, 
         -- Connections to port 'DATA11'
         DATA(10) => X_Logic0_port, 
         -- Connections to port 'DATA12'
         DATA(11) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N20, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N21, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N22, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N23, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N24, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N25, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N26, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N27, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N28, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N29, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N30, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N31, 
         -- Connections to port 'Z'
         Z(0) => N172 );
   B_0 : GTECH_BUF port map( A => N160, Z => N20);
   B_1 : GTECH_BUF port map( A => N162, Z => N21);
   B_2 : GTECH_BUF port map( A => N164, Z => N22);
   B_3 : GTECH_BUF port map( A => N166, Z => N23);
   B_4 : GTECH_BUF port map( A => N168, Z => N24);
   B_5 : GTECH_BUF port map( A => N169, Z => N25);
   B_6 : GTECH_BUF port map( A => N170, Z => N26);
   B_7 : GTECH_BUF port map( A => N171, Z => N27);
   B_8 : GTECH_BUF port map( A => N161, Z => N28);
   B_9 : GTECH_BUF port map( A => N163, Z => N29);
   B_10 : GTECH_BUF port map( A => N165, Z => N30);
   B_11 : GTECH_BUF port map( A => N167, Z => N31);
   C2007_cell : SELECT_OP
      generic map ( num_inputs => 12, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => X_Logic0_port, 
         -- Connections to port 'DATA3'
         DATA(2) => X_Logic1_port, 
         -- Connections to port 'DATA4'
         DATA(3) => X_Logic0_port, 
         -- Connections to port 'DATA5'
         DATA(4) => X_Logic1_port, 
         -- Connections to port 'DATA6'
         DATA(5) => X_Logic0_port, 
         -- Connections to port 'DATA7'
         DATA(6) => X_Logic0_port, 
         -- Connections to port 'DATA8'
         DATA(7) => X_Logic0_port, 
         -- Connections to port 'DATA9'
         DATA(8) => X_Logic1_port, 
         -- Connections to port 'DATA10'
         DATA(9) => X_Logic0_port, 
         -- Connections to port 'DATA11'
         DATA(10) => X_Logic1_port, 
         -- Connections to port 'DATA12'
         DATA(11) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N20, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N21, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N22, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N23, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N24, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N25, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N26, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N27, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N28, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N29, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N30, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N31, 
         -- Connections to port 'Z'
         Z(0) => N173 );
   C2008_cell : SELECT_OP
      generic map ( num_inputs => 12, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => X_Logic0_port, 
         -- Connections to port 'DATA3'
         DATA(2) => X_Logic1_port, 
         -- Connections to port 'DATA4'
         DATA(3) => X_Logic1_port, 
         -- Connections to port 'DATA5'
         DATA(4) => X_Logic0_port, 
         -- Connections to port 'DATA6'
         DATA(5) => X_Logic0_port, 
         -- Connections to port 'DATA7'
         DATA(6) => X_Logic0_port, 
         -- Connections to port 'DATA8'
         DATA(7) => X_Logic0_port, 
         -- Connections to port 'DATA9'
         DATA(8) => X_Logic1_port, 
         -- Connections to port 'DATA10'
         DATA(9) => X_Logic1_port, 
         -- Connections to port 'DATA11'
         DATA(10) => X_Logic1_port, 
         -- Connections to port 'DATA12'
         DATA(11) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N20, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N21, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N22, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N23, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N24, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N25, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N26, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N27, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N28, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N29, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N30, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N31, 
         -- Connections to port 'Z'
         Z(0) => N174 );
   C2009_cell : SELECT_OP
      generic map ( num_inputs => 12, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic1_port, 
         -- Connections to port 'DATA2'
         DATA(1) => X_Logic0_port, 
         -- Connections to port 'DATA3'
         DATA(2) => X_Logic1_port, 
         -- Connections to port 'DATA4'
         DATA(3) => X_Logic1_port, 
         -- Connections to port 'DATA5'
         DATA(4) => X_Logic0_port, 
         -- Connections to port 'DATA6'
         DATA(5) => X_Logic0_port, 
         -- Connections to port 'DATA7'
         DATA(6) => X_Logic1_port, 
         -- Connections to port 'DATA8'
         DATA(7) => X_Logic0_port, 
         -- Connections to port 'DATA9'
         DATA(8) => X_Logic0_port, 
         -- Connections to port 'DATA10'
         DATA(9) => X_Logic1_port, 
         -- Connections to port 'DATA11'
         DATA(10) => X_Logic0_port, 
         -- Connections to port 'DATA12'
         DATA(11) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N20, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N21, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N22, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N23, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N24, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N25, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N26, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N27, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N28, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N29, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N30, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N31, 
         -- Connections to port 'Z'
         Z(0) => N175 );
   C2010_cell : SELECT_OP
      generic map ( num_inputs => 12, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => X_Logic1_port, 
         -- Connections to port 'DATA3'
         DATA(2) => X_Logic0_port, 
         -- Connections to port 'DATA4'
         DATA(3) => X_Logic0_port, 
         -- Connections to port 'DATA5'
         DATA(4) => X_Logic1_port, 
         -- Connections to port 'DATA6'
         DATA(5) => X_Logic0_port, 
         -- Connections to port 'DATA7'
         DATA(6) => X_Logic1_port, 
         -- Connections to port 'DATA8'
         DATA(7) => X_Logic1_port, 
         -- Connections to port 'DATA9'
         DATA(8) => X_Logic0_port, 
         -- Connections to port 'DATA10'
         DATA(9) => X_Logic1_port, 
         -- Connections to port 'DATA11'
         DATA(10) => X_Logic1_port, 
         -- Connections to port 'DATA12'
         DATA(11) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N20, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N21, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N22, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N23, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N24, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N25, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N26, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N27, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N28, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N29, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N30, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N31, 
         -- Connections to port 'Z'
         Z(0) => N176 );
   C2011_cell : SELECT_OP
      generic map ( num_inputs => 12, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic1_port, 
         -- Connections to port 'DATA2'
         DATA(1) => X_Logic1_port, 
         -- Connections to port 'DATA3'
         DATA(2) => X_Logic0_port, 
         -- Connections to port 'DATA4'
         DATA(3) => X_Logic1_port, 
         -- Connections to port 'DATA5'
         DATA(4) => X_Logic0_port, 
         -- Connections to port 'DATA6'
         DATA(5) => X_Logic1_port, 
         -- Connections to port 'DATA7'
         DATA(6) => X_Logic0_port, 
         -- Connections to port 'DATA8'
         DATA(7) => X_Logic0_port, 
         -- Connections to port 'DATA9'
         DATA(8) => X_Logic0_port, 
         -- Connections to port 'DATA10'
         DATA(9) => X_Logic1_port, 
         -- Connections to port 'DATA11'
         DATA(10) => X_Logic0_port, 
         -- Connections to port 'DATA12'
         DATA(11) => X_Logic1_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N20, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N21, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N22, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N23, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N24, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N25, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N26, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N27, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N28, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N29, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N30, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N31, 
         -- Connections to port 'Z'
         Z(0) => N177 );
   C2012_cell : SELECT_OP
      generic map ( num_inputs => 12, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic1_port, 
         -- Connections to port 'DATA2'
         DATA(1) => X_Logic1_port, 
         -- Connections to port 'DATA3'
         DATA(2) => X_Logic0_port, 
         -- Connections to port 'DATA4'
         DATA(3) => X_Logic0_port, 
         -- Connections to port 'DATA5'
         DATA(4) => X_Logic0_port, 
         -- Connections to port 'DATA6'
         DATA(5) => X_Logic0_port, 
         -- Connections to port 'DATA7'
         DATA(6) => X_Logic0_port, 
         -- Connections to port 'DATA8'
         DATA(7) => X_Logic1_port, 
         -- Connections to port 'DATA9'
         DATA(8) => X_Logic0_port, 
         -- Connections to port 'DATA10'
         DATA(9) => X_Logic0_port, 
         -- Connections to port 'DATA11'
         DATA(10) => X_Logic0_port, 
         -- Connections to port 'DATA12'
         DATA(11) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N20, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N21, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N22, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N23, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N24, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N25, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N26, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N27, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N28, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N29, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N30, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N31, 
         -- Connections to port 'Z'
         Z(0) => N178 );
   C2013_cell : SELECT_OP
      generic map ( num_inputs => 12, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => X_Logic0_port, 
         -- Connections to port 'DATA3'
         DATA(2) => X_Logic0_port, 
         -- Connections to port 'DATA4'
         DATA(3) => X_Logic0_port, 
         -- Connections to port 'DATA5'
         DATA(4) => X_Logic0_port, 
         -- Connections to port 'DATA6'
         DATA(5) => X_Logic1_port, 
         -- Connections to port 'DATA7'
         DATA(6) => X_Logic0_port, 
         -- Connections to port 'DATA8'
         DATA(7) => X_Logic1_port, 
         -- Connections to port 'DATA9'
         DATA(8) => X_Logic0_port, 
         -- Connections to port 'DATA10'
         DATA(9) => X_Logic0_port, 
         -- Connections to port 'DATA11'
         DATA(10) => X_Logic0_port, 
         -- Connections to port 'DATA12'
         DATA(11) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N20, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N21, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N22, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N23, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N24, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N25, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N26, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N27, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N28, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N29, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N30, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N31, 
         -- Connections to port 'Z'
         Z(0) => N179 );
   C2014_cell : SELECT_OP
      generic map ( num_inputs => 12, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => X_Logic0_port, 
         -- Connections to port 'DATA3'
         DATA(2) => X_Logic0_port, 
         -- Connections to port 'DATA4'
         DATA(3) => X_Logic0_port, 
         -- Connections to port 'DATA5'
         DATA(4) => X_Logic0_port, 
         -- Connections to port 'DATA6'
         DATA(5) => X_Logic0_port, 
         -- Connections to port 'DATA7'
         DATA(6) => X_Logic0_port, 
         -- Connections to port 'DATA8'
         DATA(7) => X_Logic0_port, 
         -- Connections to port 'DATA9'
         DATA(8) => X_Logic0_port, 
         -- Connections to port 'DATA10'
         DATA(9) => X_Logic0_port, 
         -- Connections to port 'DATA11'
         DATA(10) => X_Logic0_port, 
         -- Connections to port 'DATA12'
         DATA(11) => X_Logic1_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N20, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N21, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N22, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N23, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N24, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N25, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N26, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N27, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N28, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N29, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N30, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N31, 
         -- Connections to port 'Z'
         Z(0) => N180 );
         X_Logic1_port <= '1';
         X_Logic0_port <= '0';
   C2017 : GTECH_XOR2 port map( A => INPUT(127), B => INPUT(255), Z => N32);
   C2018 : GTECH_XOR2 port map( A => INPUT(126), B => INPUT(254), Z => N33);
   C2019 : GTECH_XOR2 port map( A => INPUT(125), B => INPUT(253), Z => N34);
   C2020 : GTECH_XOR2 port map( A => INPUT(124), B => INPUT(252), Z => N35);
   C2021 : GTECH_XOR2 port map( A => INPUT(123), B => INPUT(251), Z => N36);
   C2022 : GTECH_XOR2 port map( A => INPUT(122), B => INPUT(250), Z => N37);
   C2023 : GTECH_XOR2 port map( A => INPUT(121), B => INPUT(249), Z => N38);
   C2024 : GTECH_XOR2 port map( A => INPUT(120), B => INPUT(248), Z => N39);
   C2025 : GTECH_XOR2 port map( A => INPUT(119), B => INPUT(247), Z => N40);
   C2026 : GTECH_XOR2 port map( A => INPUT(118), B => INPUT(246), Z => N41);
   C2027 : GTECH_XOR2 port map( A => INPUT(117), B => INPUT(245), Z => N42);
   C2028 : GTECH_XOR2 port map( A => INPUT(116), B => INPUT(244), Z => N43);
   C2029 : GTECH_XOR2 port map( A => INPUT(115), B => INPUT(243), Z => N44);
   C2030 : GTECH_XOR2 port map( A => INPUT(114), B => INPUT(242), Z => N45);
   C2031 : GTECH_XOR2 port map( A => INPUT(113), B => INPUT(241), Z => N46);
   C2032 : GTECH_XOR2 port map( A => INPUT(112), B => INPUT(240), Z => N47);
   C2033 : GTECH_XOR2 port map( A => INPUT(111), B => INPUT(239), Z => N48);
   C2034 : GTECH_XOR2 port map( A => INPUT(110), B => INPUT(238), Z => N49);
   C2035 : GTECH_XOR2 port map( A => INPUT(109), B => INPUT(237), Z => N50);
   C2036 : GTECH_XOR2 port map( A => INPUT(108), B => INPUT(236), Z => N51);
   C2037 : GTECH_XOR2 port map( A => INPUT(107), B => INPUT(235), Z => N52);
   C2038 : GTECH_XOR2 port map( A => INPUT(106), B => INPUT(234), Z => N53);
   C2039 : GTECH_XOR2 port map( A => INPUT(105), B => INPUT(233), Z => N54);
   C2040 : GTECH_XOR2 port map( A => INPUT(104), B => INPUT(232), Z => N55);
   C2041 : GTECH_XOR2 port map( A => INPUT(103), B => INPUT(231), Z => N56);
   C2042 : GTECH_XOR2 port map( A => INPUT(102), B => INPUT(230), Z => N57);
   C2043 : GTECH_XOR2 port map( A => INPUT(101), B => INPUT(229), Z => N58);
   C2044 : GTECH_XOR2 port map( A => INPUT(100), B => INPUT(228), Z => N59);
   C2045 : GTECH_XOR2 port map( A => INPUT(99), B => INPUT(227), Z => N60);
   C2046 : GTECH_XOR2 port map( A => INPUT(98), B => INPUT(226), Z => N61);
   C2047 : GTECH_XOR2 port map( A => INPUT(97), B => INPUT(225), Z => N62);
   C2048 : GTECH_XOR2 port map( A => INPUT(96), B => INPUT(224), Z => N63);
   C2049 : GTECH_XOR2 port map( A => INPUT(95), B => INPUT(223), Z => N64);
   C2050 : GTECH_XOR2 port map( A => INPUT(94), B => INPUT(222), Z => N65);
   C2051 : GTECH_XOR2 port map( A => INPUT(93), B => INPUT(221), Z => N66);
   C2052 : GTECH_XOR2 port map( A => INPUT(92), B => INPUT(220), Z => N67);
   C2053 : GTECH_XOR2 port map( A => INPUT(91), B => INPUT(219), Z => N68);
   C2054 : GTECH_XOR2 port map( A => INPUT(90), B => INPUT(218), Z => N69);
   C2055 : GTECH_XOR2 port map( A => INPUT(89), B => INPUT(217), Z => N70);
   C2056 : GTECH_XOR2 port map( A => INPUT(88), B => INPUT(216), Z => N71);
   C2057 : GTECH_XOR2 port map( A => INPUT(87), B => INPUT(215), Z => N72);
   C2058 : GTECH_XOR2 port map( A => INPUT(86), B => INPUT(214), Z => N73);
   C2059 : GTECH_XOR2 port map( A => INPUT(85), B => INPUT(213), Z => N74);
   C2060 : GTECH_XOR2 port map( A => INPUT(84), B => INPUT(212), Z => N75);
   C2061 : GTECH_XOR2 port map( A => INPUT(83), B => INPUT(211), Z => N76);
   C2062 : GTECH_XOR2 port map( A => INPUT(82), B => INPUT(210), Z => N77);
   C2063 : GTECH_XOR2 port map( A => INPUT(81), B => INPUT(209), Z => N78);
   C2064 : GTECH_XOR2 port map( A => INPUT(80), B => INPUT(208), Z => N79);
   C2065 : GTECH_XOR2 port map( A => INPUT(79), B => INPUT(207), Z => N80);
   C2066 : GTECH_XOR2 port map( A => INPUT(78), B => INPUT(206), Z => N81);
   C2067 : GTECH_XOR2 port map( A => INPUT(77), B => INPUT(205), Z => N82);
   C2068 : GTECH_XOR2 port map( A => INPUT(76), B => INPUT(204), Z => N83);
   C2069 : GTECH_XOR2 port map( A => INPUT(75), B => INPUT(203), Z => N84);
   C2070 : GTECH_XOR2 port map( A => INPUT(74), B => INPUT(202), Z => N85);
   C2071 : GTECH_XOR2 port map( A => INPUT(73), B => INPUT(201), Z => N86);
   C2072 : GTECH_XOR2 port map( A => INPUT(72), B => INPUT(200), Z => N87);
   C2073 : GTECH_XOR2 port map( A => INPUT(71), B => INPUT(199), Z => N88);
   C2074 : GTECH_XOR2 port map( A => INPUT(70), B => INPUT(198), Z => N89);
   C2075 : GTECH_XOR2 port map( A => INPUT(69), B => INPUT(197), Z => N90);
   C2076 : GTECH_XOR2 port map( A => INPUT(68), B => INPUT(196), Z => N91);
   C2077 : GTECH_XOR2 port map( A => INPUT(67), B => INPUT(195), Z => N92);
   C2078 : GTECH_XOR2 port map( A => INPUT(66), B => INPUT(194), Z => N93);
   C2079 : GTECH_XOR2 port map( A => INPUT(65), B => INPUT(193), Z => N94);
   C2080 : GTECH_XOR2 port map( A => INPUT(64), B => INPUT(192), Z => N95);
   C2081 : GTECH_XOR2 port map( A => INPUT(63), B => INPUT(191), Z => N96);
   C2082 : GTECH_XOR2 port map( A => INPUT(62), B => INPUT(190), Z => N97);
   C2083 : GTECH_XOR2 port map( A => INPUT(61), B => INPUT(189), Z => N98);
   C2084 : GTECH_XOR2 port map( A => INPUT(60), B => INPUT(188), Z => N99);
   C2085 : GTECH_XOR2 port map( A => INPUT(59), B => INPUT(187), Z => N100);
   C2086 : GTECH_XOR2 port map( A => INPUT(58), B => INPUT(186), Z => N101);
   C2087 : GTECH_XOR2 port map( A => INPUT(57), B => INPUT(185), Z => N102);
   C2088 : GTECH_XOR2 port map( A => INPUT(56), B => INPUT(184), Z => N103);
   C2089 : GTECH_XOR2 port map( A => INPUT(55), B => INPUT(183), Z => N104);
   C2090 : GTECH_XOR2 port map( A => INPUT(54), B => INPUT(182), Z => N105);
   C2091 : GTECH_XOR2 port map( A => INPUT(53), B => INPUT(181), Z => N106);
   C2092 : GTECH_XOR2 port map( A => INPUT(52), B => INPUT(180), Z => N107);
   C2093 : GTECH_XOR2 port map( A => INPUT(51), B => INPUT(179), Z => N108);
   C2094 : GTECH_XOR2 port map( A => INPUT(50), B => INPUT(178), Z => N109);
   C2095 : GTECH_XOR2 port map( A => INPUT(49), B => INPUT(177), Z => N110);
   C2096 : GTECH_XOR2 port map( A => INPUT(48), B => INPUT(176), Z => N111);
   C2097 : GTECH_XOR2 port map( A => INPUT(47), B => INPUT(175), Z => N112);
   C2098 : GTECH_XOR2 port map( A => INPUT(46), B => INPUT(174), Z => N113);
   C2099 : GTECH_XOR2 port map( A => INPUT(45), B => INPUT(173), Z => N114);
   C2100 : GTECH_XOR2 port map( A => INPUT(44), B => INPUT(172), Z => N115);
   C2101 : GTECH_XOR2 port map( A => INPUT(43), B => INPUT(171), Z => N116);
   C2102 : GTECH_XOR2 port map( A => INPUT(42), B => INPUT(170), Z => N117);
   C2103 : GTECH_XOR2 port map( A => INPUT(41), B => INPUT(169), Z => N118);
   C2104 : GTECH_XOR2 port map( A => INPUT(40), B => INPUT(168), Z => N119);
   C2105 : GTECH_XOR2 port map( A => INPUT(39), B => INPUT(167), Z => N120);
   C2106 : GTECH_XOR2 port map( A => INPUT(38), B => INPUT(166), Z => N121);
   C2107 : GTECH_XOR2 port map( A => INPUT(37), B => INPUT(165), Z => N122);
   C2108 : GTECH_XOR2 port map( A => INPUT(36), B => INPUT(164), Z => N123);
   C2109 : GTECH_XOR2 port map( A => INPUT(35), B => INPUT(163), Z => N124);
   C2110 : GTECH_XOR2 port map( A => INPUT(34), B => INPUT(162), Z => N125);
   C2111 : GTECH_XOR2 port map( A => INPUT(33), B => INPUT(161), Z => N126);
   C2112 : GTECH_XOR2 port map( A => INPUT(32), B => INPUT(160), Z => N127);
   C2113 : GTECH_XOR2 port map( A => INPUT(31), B => INPUT(159), Z => N128);
   C2114 : GTECH_XOR2 port map( A => INPUT(30), B => INPUT(158), Z => N129);
   C2115 : GTECH_XOR2 port map( A => INPUT(29), B => INPUT(157), Z => N130);
   C2116 : GTECH_XOR2 port map( A => INPUT(28), B => INPUT(156), Z => N131);
   C2117 : GTECH_XOR2 port map( A => INPUT(27), B => INPUT(155), Z => N132);
   C2118 : GTECH_XOR2 port map( A => INPUT(26), B => INPUT(154), Z => N133);
   C2119 : GTECH_XOR2 port map( A => INPUT(25), B => INPUT(153), Z => N134);
   C2120 : GTECH_XOR2 port map( A => INPUT(24), B => INPUT(152), Z => N135);
   C2121 : GTECH_XOR2 port map( A => INPUT(23), B => INPUT(151), Z => N136);
   C2122 : GTECH_XOR2 port map( A => INPUT(22), B => INPUT(150), Z => N137);
   C2123 : GTECH_XOR2 port map( A => INPUT(21), B => INPUT(149), Z => N138);
   C2124 : GTECH_XOR2 port map( A => INPUT(20), B => INPUT(148), Z => N139);
   C2125 : GTECH_XOR2 port map( A => INPUT(19), B => INPUT(147), Z => N140);
   C2126 : GTECH_XOR2 port map( A => INPUT(18), B => INPUT(146), Z => N141);
   C2127 : GTECH_XOR2 port map( A => INPUT(17), B => INPUT(145), Z => N142);
   C2128 : GTECH_XOR2 port map( A => INPUT(16), B => INPUT(144), Z => N143);
   C2129 : GTECH_XOR2 port map( A => INPUT(15), B => INPUT(143), Z => N144);
   C2130 : GTECH_XOR2 port map( A => INPUT(14), B => INPUT(142), Z => N145);
   C2131 : GTECH_XOR2 port map( A => INPUT(13), B => INPUT(141), Z => N146);
   C2132 : GTECH_XOR2 port map( A => INPUT(12), B => INPUT(140), Z => N147);
   C2133 : GTECH_XOR2 port map( A => INPUT(11), B => INPUT(139), Z => N148);
   C2134 : GTECH_XOR2 port map( A => INPUT(10), B => INPUT(138), Z => N149);
   C2135 : GTECH_XOR2 port map( A => INPUT(9), B => INPUT(137), Z => N150);
   C2136 : GTECH_XOR2 port map( A => INPUT(8), B => INPUT(136), Z => N151);
   C2137 : GTECH_XOR2 port map( A => INPUT(7), B => INPUT(135), Z => N152);
   C2138 : GTECH_XOR2 port map( A => INPUT(6), B => INPUT(134), Z => N153);
   C2139 : GTECH_XOR2 port map( A => INPUT(5), B => INPUT(133), Z => N154);
   C2140 : GTECH_XOR2 port map( A => INPUT(4), B => INPUT(132), Z => N155);
   C2141 : GTECH_XOR2 port map( A => INPUT(3), B => INPUT(131), Z => N156);
   C2142 : GTECH_XOR2 port map( A => INPUT(2), B => INPUT(130), Z => N157);
   C2143 : GTECH_XOR2 port map( A => INPUT(1), B => INPUT(129), Z => N158);
   C2144 : GTECH_XOR2 port map( A => INPUT(0), B => INPUT(128), Z => N159);
   C2145 : GTECH_XOR2 port map( A => N32, B => INPUT(383), Z => 
                           p_plane_127_port);
   C2146 : GTECH_XOR2 port map( A => N33, B => INPUT(382), Z => 
                           p_plane_126_port);
   C2147 : GTECH_XOR2 port map( A => N34, B => INPUT(381), Z => 
                           p_plane_125_port);
   C2148 : GTECH_XOR2 port map( A => N35, B => INPUT(380), Z => 
                           p_plane_124_port);
   C2149 : GTECH_XOR2 port map( A => N36, B => INPUT(379), Z => 
                           p_plane_123_port);
   C2150 : GTECH_XOR2 port map( A => N37, B => INPUT(378), Z => 
                           p_plane_122_port);
   C2151 : GTECH_XOR2 port map( A => N38, B => INPUT(377), Z => 
                           p_plane_121_port);
   C2152 : GTECH_XOR2 port map( A => N39, B => INPUT(376), Z => 
                           p_plane_120_port);
   C2153 : GTECH_XOR2 port map( A => N40, B => INPUT(375), Z => 
                           p_plane_119_port);
   C2154 : GTECH_XOR2 port map( A => N41, B => INPUT(374), Z => 
                           p_plane_118_port);
   C2155 : GTECH_XOR2 port map( A => N42, B => INPUT(373), Z => 
                           p_plane_117_port);
   C2156 : GTECH_XOR2 port map( A => N43, B => INPUT(372), Z => 
                           p_plane_116_port);
   C2157 : GTECH_XOR2 port map( A => N44, B => INPUT(371), Z => 
                           p_plane_115_port);
   C2158 : GTECH_XOR2 port map( A => N45, B => INPUT(370), Z => 
                           p_plane_114_port);
   C2159 : GTECH_XOR2 port map( A => N46, B => INPUT(369), Z => 
                           p_plane_113_port);
   C2160 : GTECH_XOR2 port map( A => N47, B => INPUT(368), Z => 
                           p_plane_112_port);
   C2161 : GTECH_XOR2 port map( A => N48, B => INPUT(367), Z => 
                           p_plane_111_port);
   C2162 : GTECH_XOR2 port map( A => N49, B => INPUT(366), Z => 
                           p_plane_110_port);
   C2163 : GTECH_XOR2 port map( A => N50, B => INPUT(365), Z => 
                           p_plane_109_port);
   C2164 : GTECH_XOR2 port map( A => N51, B => INPUT(364), Z => 
                           p_plane_108_port);
   C2165 : GTECH_XOR2 port map( A => N52, B => INPUT(363), Z => 
                           p_plane_107_port);
   C2166 : GTECH_XOR2 port map( A => N53, B => INPUT(362), Z => 
                           p_plane_106_port);
   C2167 : GTECH_XOR2 port map( A => N54, B => INPUT(361), Z => 
                           p_plane_105_port);
   C2168 : GTECH_XOR2 port map( A => N55, B => INPUT(360), Z => 
                           p_plane_104_port);
   C2169 : GTECH_XOR2 port map( A => N56, B => INPUT(359), Z => 
                           p_plane_103_port);
   C2170 : GTECH_XOR2 port map( A => N57, B => INPUT(358), Z => 
                           p_plane_102_port);
   C2171 : GTECH_XOR2 port map( A => N58, B => INPUT(357), Z => 
                           p_plane_101_port);
   C2172 : GTECH_XOR2 port map( A => N59, B => INPUT(356), Z => 
                           p_plane_100_port);
   C2173 : GTECH_XOR2 port map( A => N60, B => INPUT(355), Z => p_plane_99_port
                           );
   C2174 : GTECH_XOR2 port map( A => N61, B => INPUT(354), Z => p_plane_98_port
                           );
   C2175 : GTECH_XOR2 port map( A => N62, B => INPUT(353), Z => p_plane_97_port
                           );
   C2176 : GTECH_XOR2 port map( A => N63, B => INPUT(352), Z => p_plane_96_port
                           );
   C2177 : GTECH_XOR2 port map( A => N64, B => INPUT(351), Z => p_plane_95_port
                           );
   C2178 : GTECH_XOR2 port map( A => N65, B => INPUT(350), Z => p_plane_94_port
                           );
   C2179 : GTECH_XOR2 port map( A => N66, B => INPUT(349), Z => p_plane_93_port
                           );
   C2180 : GTECH_XOR2 port map( A => N67, B => INPUT(348), Z => p_plane_92_port
                           );
   C2181 : GTECH_XOR2 port map( A => N68, B => INPUT(347), Z => p_plane_91_port
                           );
   C2182 : GTECH_XOR2 port map( A => N69, B => INPUT(346), Z => p_plane_90_port
                           );
   C2183 : GTECH_XOR2 port map( A => N70, B => INPUT(345), Z => p_plane_89_port
                           );
   C2184 : GTECH_XOR2 port map( A => N71, B => INPUT(344), Z => p_plane_88_port
                           );
   C2185 : GTECH_XOR2 port map( A => N72, B => INPUT(343), Z => p_plane_87_port
                           );
   C2186 : GTECH_XOR2 port map( A => N73, B => INPUT(342), Z => p_plane_86_port
                           );
   C2187 : GTECH_XOR2 port map( A => N74, B => INPUT(341), Z => p_plane_85_port
                           );
   C2188 : GTECH_XOR2 port map( A => N75, B => INPUT(340), Z => p_plane_84_port
                           );
   C2189 : GTECH_XOR2 port map( A => N76, B => INPUT(339), Z => p_plane_83_port
                           );
   C2190 : GTECH_XOR2 port map( A => N77, B => INPUT(338), Z => p_plane_82_port
                           );
   C2191 : GTECH_XOR2 port map( A => N78, B => INPUT(337), Z => p_plane_81_port
                           );
   C2192 : GTECH_XOR2 port map( A => N79, B => INPUT(336), Z => p_plane_80_port
                           );
   C2193 : GTECH_XOR2 port map( A => N80, B => INPUT(335), Z => p_plane_79_port
                           );
   C2194 : GTECH_XOR2 port map( A => N81, B => INPUT(334), Z => p_plane_78_port
                           );
   C2195 : GTECH_XOR2 port map( A => N82, B => INPUT(333), Z => p_plane_77_port
                           );
   C2196 : GTECH_XOR2 port map( A => N83, B => INPUT(332), Z => p_plane_76_port
                           );
   C2197 : GTECH_XOR2 port map( A => N84, B => INPUT(331), Z => p_plane_75_port
                           );
   C2198 : GTECH_XOR2 port map( A => N85, B => INPUT(330), Z => p_plane_74_port
                           );
   C2199 : GTECH_XOR2 port map( A => N86, B => INPUT(329), Z => p_plane_73_port
                           );
   C2200 : GTECH_XOR2 port map( A => N87, B => INPUT(328), Z => p_plane_72_port
                           );
   C2201 : GTECH_XOR2 port map( A => N88, B => INPUT(327), Z => p_plane_71_port
                           );
   C2202 : GTECH_XOR2 port map( A => N89, B => INPUT(326), Z => p_plane_70_port
                           );
   C2203 : GTECH_XOR2 port map( A => N90, B => INPUT(325), Z => p_plane_69_port
                           );
   C2204 : GTECH_XOR2 port map( A => N91, B => INPUT(324), Z => p_plane_68_port
                           );
   C2205 : GTECH_XOR2 port map( A => N92, B => INPUT(323), Z => p_plane_67_port
                           );
   C2206 : GTECH_XOR2 port map( A => N93, B => INPUT(322), Z => p_plane_66_port
                           );
   C2207 : GTECH_XOR2 port map( A => N94, B => INPUT(321), Z => p_plane_65_port
                           );
   C2208 : GTECH_XOR2 port map( A => N95, B => INPUT(320), Z => p_plane_64_port
                           );
   C2209 : GTECH_XOR2 port map( A => N96, B => INPUT(319), Z => p_plane_63_port
                           );
   C2210 : GTECH_XOR2 port map( A => N97, B => INPUT(318), Z => p_plane_62_port
                           );
   C2211 : GTECH_XOR2 port map( A => N98, B => INPUT(317), Z => p_plane_61_port
                           );
   C2212 : GTECH_XOR2 port map( A => N99, B => INPUT(316), Z => p_plane_60_port
                           );
   C2213 : GTECH_XOR2 port map( A => N100, B => INPUT(315), Z => 
                           p_plane_59_port);
   C2214 : GTECH_XOR2 port map( A => N101, B => INPUT(314), Z => 
                           p_plane_58_port);
   C2215 : GTECH_XOR2 port map( A => N102, B => INPUT(313), Z => 
                           p_plane_57_port);
   C2216 : GTECH_XOR2 port map( A => N103, B => INPUT(312), Z => 
                           p_plane_56_port);
   C2217 : GTECH_XOR2 port map( A => N104, B => INPUT(311), Z => 
                           p_plane_55_port);
   C2218 : GTECH_XOR2 port map( A => N105, B => INPUT(310), Z => 
                           p_plane_54_port);
   C2219 : GTECH_XOR2 port map( A => N106, B => INPUT(309), Z => 
                           p_plane_53_port);
   C2220 : GTECH_XOR2 port map( A => N107, B => INPUT(308), Z => 
                           p_plane_52_port);
   C2221 : GTECH_XOR2 port map( A => N108, B => INPUT(307), Z => 
                           p_plane_51_port);
   C2222 : GTECH_XOR2 port map( A => N109, B => INPUT(306), Z => 
                           p_plane_50_port);
   C2223 : GTECH_XOR2 port map( A => N110, B => INPUT(305), Z => 
                           p_plane_49_port);
   C2224 : GTECH_XOR2 port map( A => N111, B => INPUT(304), Z => 
                           p_plane_48_port);
   C2225 : GTECH_XOR2 port map( A => N112, B => INPUT(303), Z => 
                           p_plane_47_port);
   C2226 : GTECH_XOR2 port map( A => N113, B => INPUT(302), Z => 
                           p_plane_46_port);
   C2227 : GTECH_XOR2 port map( A => N114, B => INPUT(301), Z => 
                           p_plane_45_port);
   C2228 : GTECH_XOR2 port map( A => N115, B => INPUT(300), Z => 
                           p_plane_44_port);
   C2229 : GTECH_XOR2 port map( A => N116, B => INPUT(299), Z => 
                           p_plane_43_port);
   C2230 : GTECH_XOR2 port map( A => N117, B => INPUT(298), Z => 
                           p_plane_42_port);
   C2231 : GTECH_XOR2 port map( A => N118, B => INPUT(297), Z => 
                           p_plane_41_port);
   C2232 : GTECH_XOR2 port map( A => N119, B => INPUT(296), Z => 
                           p_plane_40_port);
   C2233 : GTECH_XOR2 port map( A => N120, B => INPUT(295), Z => 
                           p_plane_39_port);
   C2234 : GTECH_XOR2 port map( A => N121, B => INPUT(294), Z => 
                           p_plane_38_port);
   C2235 : GTECH_XOR2 port map( A => N122, B => INPUT(293), Z => 
                           p_plane_37_port);
   C2236 : GTECH_XOR2 port map( A => N123, B => INPUT(292), Z => 
                           p_plane_36_port);
   C2237 : GTECH_XOR2 port map( A => N124, B => INPUT(291), Z => 
                           p_plane_35_port);
   C2238 : GTECH_XOR2 port map( A => N125, B => INPUT(290), Z => 
                           p_plane_34_port);
   C2239 : GTECH_XOR2 port map( A => N126, B => INPUT(289), Z => 
                           p_plane_33_port);
   C2240 : GTECH_XOR2 port map( A => N127, B => INPUT(288), Z => 
                           p_plane_32_port);
   C2241 : GTECH_XOR2 port map( A => N128, B => INPUT(287), Z => 
                           p_plane_31_port);
   C2242 : GTECH_XOR2 port map( A => N129, B => INPUT(286), Z => 
                           p_plane_30_port);
   C2243 : GTECH_XOR2 port map( A => N130, B => INPUT(285), Z => 
                           p_plane_29_port);
   C2244 : GTECH_XOR2 port map( A => N131, B => INPUT(284), Z => 
                           p_plane_28_port);
   C2245 : GTECH_XOR2 port map( A => N132, B => INPUT(283), Z => 
                           p_plane_27_port);
   C2246 : GTECH_XOR2 port map( A => N133, B => INPUT(282), Z => 
                           p_plane_26_port);
   C2247 : GTECH_XOR2 port map( A => N134, B => INPUT(281), Z => 
                           p_plane_25_port);
   C2248 : GTECH_XOR2 port map( A => N135, B => INPUT(280), Z => 
                           p_plane_24_port);
   C2249 : GTECH_XOR2 port map( A => N136, B => INPUT(279), Z => 
                           p_plane_23_port);
   C2250 : GTECH_XOR2 port map( A => N137, B => INPUT(278), Z => 
                           p_plane_22_port);
   C2251 : GTECH_XOR2 port map( A => N138, B => INPUT(277), Z => 
                           p_plane_21_port);
   C2252 : GTECH_XOR2 port map( A => N139, B => INPUT(276), Z => 
                           p_plane_20_port);
   C2253 : GTECH_XOR2 port map( A => N140, B => INPUT(275), Z => 
                           p_plane_19_port);
   C2254 : GTECH_XOR2 port map( A => N141, B => INPUT(274), Z => 
                           p_plane_18_port);
   C2255 : GTECH_XOR2 port map( A => N142, B => INPUT(273), Z => 
                           p_plane_17_port);
   C2256 : GTECH_XOR2 port map( A => N143, B => INPUT(272), Z => 
                           p_plane_16_port);
   C2257 : GTECH_XOR2 port map( A => N144, B => INPUT(271), Z => 
                           p_plane_15_port);
   C2258 : GTECH_XOR2 port map( A => N145, B => INPUT(270), Z => 
                           p_plane_14_port);
   C2259 : GTECH_XOR2 port map( A => N146, B => INPUT(269), Z => 
                           p_plane_13_port);
   C2260 : GTECH_XOR2 port map( A => N147, B => INPUT(268), Z => 
                           p_plane_12_port);
   C2261 : GTECH_XOR2 port map( A => N148, B => INPUT(267), Z => 
                           p_plane_11_port);
   C2262 : GTECH_XOR2 port map( A => N149, B => INPUT(266), Z => 
                           p_plane_10_port);
   C2263 : GTECH_XOR2 port map( A => N150, B => INPUT(265), Z => p_plane_9_port
                           );
   C2264 : GTECH_XOR2 port map( A => N151, B => INPUT(264), Z => p_plane_8_port
                           );
   C2265 : GTECH_XOR2 port map( A => N152, B => INPUT(263), Z => p_plane_7_port
                           );
   C2266 : GTECH_XOR2 port map( A => N153, B => INPUT(262), Z => p_plane_6_port
                           );
   C2267 : GTECH_XOR2 port map( A => N154, B => INPUT(261), Z => p_plane_5_port
                           );
   C2268 : GTECH_XOR2 port map( A => N155, B => INPUT(260), Z => p_plane_4_port
                           );
   C2269 : GTECH_XOR2 port map( A => N156, B => INPUT(259), Z => p_plane_3_port
                           );
   C2270 : GTECH_XOR2 port map( A => N157, B => INPUT(258), Z => p_plane_2_port
                           );
   C2271 : GTECH_XOR2 port map( A => N158, B => INPUT(257), Z => p_plane_1_port
                           );
   C2272 : GTECH_XOR2 port map( A => N159, B => INPUT(256), Z => p_plane_0_port
                           );
   C2273 : GTECH_XOR2 port map( A => p_plane_26_port, B => p_plane_17_port, Z 
                           => eshift_127_port);
   C2274 : GTECH_XOR2 port map( A => p_plane_25_port, B => p_plane_16_port, Z 
                           => eshift_126_port);
   C2275 : GTECH_XOR2 port map( A => p_plane_24_port, B => p_plane_15_port, Z 
                           => eshift_125_port);
   C2276 : GTECH_XOR2 port map( A => p_plane_23_port, B => p_plane_14_port, Z 
                           => eshift_124_port);
   C2277 : GTECH_XOR2 port map( A => p_plane_22_port, B => p_plane_13_port, Z 
                           => eshift_123_port);
   C2278 : GTECH_XOR2 port map( A => p_plane_21_port, B => p_plane_12_port, Z 
                           => eshift_122_port);
   C2279 : GTECH_XOR2 port map( A => p_plane_20_port, B => p_plane_11_port, Z 
                           => eshift_121_port);
   C2280 : GTECH_XOR2 port map( A => p_plane_19_port, B => p_plane_10_port, Z 
                           => eshift_120_port);
   C2281 : GTECH_XOR2 port map( A => p_plane_18_port, B => p_plane_9_port, Z =>
                           eshift_119_port);
   C2282 : GTECH_XOR2 port map( A => p_plane_17_port, B => p_plane_8_port, Z =>
                           eshift_118_port);
   C2283 : GTECH_XOR2 port map( A => p_plane_16_port, B => p_plane_7_port, Z =>
                           eshift_117_port);
   C2284 : GTECH_XOR2 port map( A => p_plane_15_port, B => p_plane_6_port, Z =>
                           eshift_116_port);
   C2285 : GTECH_XOR2 port map( A => p_plane_14_port, B => p_plane_5_port, Z =>
                           eshift_115_port);
   C2286 : GTECH_XOR2 port map( A => p_plane_13_port, B => p_plane_4_port, Z =>
                           eshift_114_port);
   C2287 : GTECH_XOR2 port map( A => p_plane_12_port, B => p_plane_3_port, Z =>
                           eshift_113_port);
   C2288 : GTECH_XOR2 port map( A => p_plane_11_port, B => p_plane_2_port, Z =>
                           eshift_112_port);
   C2289 : GTECH_XOR2 port map( A => p_plane_10_port, B => p_plane_1_port, Z =>
                           eshift_111_port);
   C2290 : GTECH_XOR2 port map( A => p_plane_9_port, B => p_plane_0_port, Z => 
                           eshift_110_port);
   C2291 : GTECH_XOR2 port map( A => p_plane_8_port, B => p_plane_31_port, Z =>
                           eshift_109_port);
   C2292 : GTECH_XOR2 port map( A => p_plane_7_port, B => p_plane_30_port, Z =>
                           eshift_108_port);
   C2293 : GTECH_XOR2 port map( A => p_plane_6_port, B => p_plane_29_port, Z =>
                           eshift_107_port);
   C2294 : GTECH_XOR2 port map( A => p_plane_5_port, B => p_plane_28_port, Z =>
                           eshift_106_port);
   C2295 : GTECH_XOR2 port map( A => p_plane_4_port, B => p_plane_27_port, Z =>
                           eshift_105_port);
   C2296 : GTECH_XOR2 port map( A => p_plane_3_port, B => p_plane_26_port, Z =>
                           eshift_104_port);
   C2297 : GTECH_XOR2 port map( A => p_plane_2_port, B => p_plane_25_port, Z =>
                           eshift_103_port);
   C2298 : GTECH_XOR2 port map( A => p_plane_1_port, B => p_plane_24_port, Z =>
                           eshift_102_port);
   C2299 : GTECH_XOR2 port map( A => p_plane_0_port, B => p_plane_23_port, Z =>
                           eshift_101_port);
   C2300 : GTECH_XOR2 port map( A => p_plane_31_port, B => p_plane_22_port, Z 
                           => eshift_100_port);
   C2301 : GTECH_XOR2 port map( A => p_plane_30_port, B => p_plane_21_port, Z 
                           => eshift_99_port);
   C2302 : GTECH_XOR2 port map( A => p_plane_29_port, B => p_plane_20_port, Z 
                           => eshift_98_port);
   C2303 : GTECH_XOR2 port map( A => p_plane_28_port, B => p_plane_19_port, Z 
                           => eshift_97_port);
   C2304 : GTECH_XOR2 port map( A => p_plane_27_port, B => p_plane_18_port, Z 
                           => eshift_96_port);
   C2305 : GTECH_XOR2 port map( A => p_plane_122_port, B => p_plane_113_port, Z
                           => eshift_95_port);
   C2306 : GTECH_XOR2 port map( A => p_plane_121_port, B => p_plane_112_port, Z
                           => eshift_94_port);
   C2307 : GTECH_XOR2 port map( A => p_plane_120_port, B => p_plane_111_port, Z
                           => eshift_93_port);
   C2308 : GTECH_XOR2 port map( A => p_plane_119_port, B => p_plane_110_port, Z
                           => eshift_92_port);
   C2309 : GTECH_XOR2 port map( A => p_plane_118_port, B => p_plane_109_port, Z
                           => eshift_91_port);
   C2310 : GTECH_XOR2 port map( A => p_plane_117_port, B => p_plane_108_port, Z
                           => eshift_90_port);
   C2311 : GTECH_XOR2 port map( A => p_plane_116_port, B => p_plane_107_port, Z
                           => eshift_89_port);
   C2312 : GTECH_XOR2 port map( A => p_plane_115_port, B => p_plane_106_port, Z
                           => eshift_88_port);
   C2313 : GTECH_XOR2 port map( A => p_plane_114_port, B => p_plane_105_port, Z
                           => eshift_87_port);
   C2314 : GTECH_XOR2 port map( A => p_plane_113_port, B => p_plane_104_port, Z
                           => eshift_86_port);
   C2315 : GTECH_XOR2 port map( A => p_plane_112_port, B => p_plane_103_port, Z
                           => eshift_85_port);
   C2316 : GTECH_XOR2 port map( A => p_plane_111_port, B => p_plane_102_port, Z
                           => eshift_84_port);
   C2317 : GTECH_XOR2 port map( A => p_plane_110_port, B => p_plane_101_port, Z
                           => eshift_83_port);
   C2318 : GTECH_XOR2 port map( A => p_plane_109_port, B => p_plane_100_port, Z
                           => eshift_82_port);
   C2319 : GTECH_XOR2 port map( A => p_plane_108_port, B => p_plane_99_port, Z 
                           => eshift_81_port);
   C2320 : GTECH_XOR2 port map( A => p_plane_107_port, B => p_plane_98_port, Z 
                           => eshift_80_port);
   C2321 : GTECH_XOR2 port map( A => p_plane_106_port, B => p_plane_97_port, Z 
                           => eshift_79_port);
   C2322 : GTECH_XOR2 port map( A => p_plane_105_port, B => p_plane_96_port, Z 
                           => eshift_78_port);
   C2323 : GTECH_XOR2 port map( A => p_plane_104_port, B => p_plane_127_port, Z
                           => eshift_77_port);
   C2324 : GTECH_XOR2 port map( A => p_plane_103_port, B => p_plane_126_port, Z
                           => eshift_76_port);
   C2325 : GTECH_XOR2 port map( A => p_plane_102_port, B => p_plane_125_port, Z
                           => eshift_75_port);
   C2326 : GTECH_XOR2 port map( A => p_plane_101_port, B => p_plane_124_port, Z
                           => eshift_74_port);
   C2327 : GTECH_XOR2 port map( A => p_plane_100_port, B => p_plane_123_port, Z
                           => eshift_73_port);
   C2328 : GTECH_XOR2 port map( A => p_plane_99_port, B => p_plane_122_port, Z 
                           => eshift_72_port);
   C2329 : GTECH_XOR2 port map( A => p_plane_98_port, B => p_plane_121_port, Z 
                           => eshift_71_port);
   C2330 : GTECH_XOR2 port map( A => p_plane_97_port, B => p_plane_120_port, Z 
                           => eshift_70_port);
   C2331 : GTECH_XOR2 port map( A => p_plane_96_port, B => p_plane_119_port, Z 
                           => eshift_69_port);
   C2332 : GTECH_XOR2 port map( A => p_plane_127_port, B => p_plane_118_port, Z
                           => eshift_68_port);
   C2333 : GTECH_XOR2 port map( A => p_plane_126_port, B => p_plane_117_port, Z
                           => eshift_67_port);
   C2334 : GTECH_XOR2 port map( A => p_plane_125_port, B => p_plane_116_port, Z
                           => eshift_66_port);
   C2335 : GTECH_XOR2 port map( A => p_plane_124_port, B => p_plane_115_port, Z
                           => eshift_65_port);
   C2336 : GTECH_XOR2 port map( A => p_plane_123_port, B => p_plane_114_port, Z
                           => eshift_64_port);
   C2337 : GTECH_XOR2 port map( A => p_plane_90_port, B => p_plane_81_port, Z 
                           => eshift_63_port);
   C2338 : GTECH_XOR2 port map( A => p_plane_89_port, B => p_plane_80_port, Z 
                           => eshift_62_port);
   C2339 : GTECH_XOR2 port map( A => p_plane_88_port, B => p_plane_79_port, Z 
                           => eshift_61_port);
   C2340 : GTECH_XOR2 port map( A => p_plane_87_port, B => p_plane_78_port, Z 
                           => eshift_60_port);
   C2341 : GTECH_XOR2 port map( A => p_plane_86_port, B => p_plane_77_port, Z 
                           => eshift_59_port);
   C2342 : GTECH_XOR2 port map( A => p_plane_85_port, B => p_plane_76_port, Z 
                           => eshift_58_port);
   C2343 : GTECH_XOR2 port map( A => p_plane_84_port, B => p_plane_75_port, Z 
                           => eshift_57_port);
   C2344 : GTECH_XOR2 port map( A => p_plane_83_port, B => p_plane_74_port, Z 
                           => eshift_56_port);
   C2345 : GTECH_XOR2 port map( A => p_plane_82_port, B => p_plane_73_port, Z 
                           => eshift_55_port);
   C2346 : GTECH_XOR2 port map( A => p_plane_81_port, B => p_plane_72_port, Z 
                           => eshift_54_port);
   C2347 : GTECH_XOR2 port map( A => p_plane_80_port, B => p_plane_71_port, Z 
                           => eshift_53_port);
   C2348 : GTECH_XOR2 port map( A => p_plane_79_port, B => p_plane_70_port, Z 
                           => eshift_52_port);
   C2349 : GTECH_XOR2 port map( A => p_plane_78_port, B => p_plane_69_port, Z 
                           => eshift_51_port);
   C2350 : GTECH_XOR2 port map( A => p_plane_77_port, B => p_plane_68_port, Z 
                           => eshift_50_port);
   C2351 : GTECH_XOR2 port map( A => p_plane_76_port, B => p_plane_67_port, Z 
                           => eshift_49_port);
   C2352 : GTECH_XOR2 port map( A => p_plane_75_port, B => p_plane_66_port, Z 
                           => eshift_48_port);
   C2353 : GTECH_XOR2 port map( A => p_plane_74_port, B => p_plane_65_port, Z 
                           => eshift_47_port);
   C2354 : GTECH_XOR2 port map( A => p_plane_73_port, B => p_plane_64_port, Z 
                           => eshift_46_port);
   C2355 : GTECH_XOR2 port map( A => p_plane_72_port, B => p_plane_95_port, Z 
                           => eshift_45_port);
   C2356 : GTECH_XOR2 port map( A => p_plane_71_port, B => p_plane_94_port, Z 
                           => eshift_44_port);
   C2357 : GTECH_XOR2 port map( A => p_plane_70_port, B => p_plane_93_port, Z 
                           => eshift_43_port);
   C2358 : GTECH_XOR2 port map( A => p_plane_69_port, B => p_plane_92_port, Z 
                           => eshift_42_port);
   C2359 : GTECH_XOR2 port map( A => p_plane_68_port, B => p_plane_91_port, Z 
                           => eshift_41_port);
   C2360 : GTECH_XOR2 port map( A => p_plane_67_port, B => p_plane_90_port, Z 
                           => eshift_40_port);
   C2361 : GTECH_XOR2 port map( A => p_plane_66_port, B => p_plane_89_port, Z 
                           => eshift_39_port);
   C2362 : GTECH_XOR2 port map( A => p_plane_65_port, B => p_plane_88_port, Z 
                           => eshift_38_port);
   C2363 : GTECH_XOR2 port map( A => p_plane_64_port, B => p_plane_87_port, Z 
                           => eshift_37_port);
   C2364 : GTECH_XOR2 port map( A => p_plane_95_port, B => p_plane_86_port, Z 
                           => eshift_36_port);
   C2365 : GTECH_XOR2 port map( A => p_plane_94_port, B => p_plane_85_port, Z 
                           => eshift_35_port);
   C2366 : GTECH_XOR2 port map( A => p_plane_93_port, B => p_plane_84_port, Z 
                           => eshift_34_port);
   C2367 : GTECH_XOR2 port map( A => p_plane_92_port, B => p_plane_83_port, Z 
                           => eshift_33_port);
   C2368 : GTECH_XOR2 port map( A => p_plane_91_port, B => p_plane_82_port, Z 
                           => eshift_32_port);
   C2369 : GTECH_XOR2 port map( A => p_plane_58_port, B => p_plane_49_port, Z 
                           => eshift_31_port);
   C2370 : GTECH_XOR2 port map( A => p_plane_57_port, B => p_plane_48_port, Z 
                           => eshift_30_port);
   C2371 : GTECH_XOR2 port map( A => p_plane_56_port, B => p_plane_47_port, Z 
                           => eshift_29_port);
   C2372 : GTECH_XOR2 port map( A => p_plane_55_port, B => p_plane_46_port, Z 
                           => eshift_28_port);
   C2373 : GTECH_XOR2 port map( A => p_plane_54_port, B => p_plane_45_port, Z 
                           => eshift_27_port);
   C2374 : GTECH_XOR2 port map( A => p_plane_53_port, B => p_plane_44_port, Z 
                           => eshift_26_port);
   C2375 : GTECH_XOR2 port map( A => p_plane_52_port, B => p_plane_43_port, Z 
                           => eshift_25_port);
   C2376 : GTECH_XOR2 port map( A => p_plane_51_port, B => p_plane_42_port, Z 
                           => eshift_24_port);
   C2377 : GTECH_XOR2 port map( A => p_plane_50_port, B => p_plane_41_port, Z 
                           => eshift_23_port);
   C2378 : GTECH_XOR2 port map( A => p_plane_49_port, B => p_plane_40_port, Z 
                           => eshift_22_port);
   C2379 : GTECH_XOR2 port map( A => p_plane_48_port, B => p_plane_39_port, Z 
                           => eshift_21_port);
   C2380 : GTECH_XOR2 port map( A => p_plane_47_port, B => p_plane_38_port, Z 
                           => eshift_20_port);
   C2381 : GTECH_XOR2 port map( A => p_plane_46_port, B => p_plane_37_port, Z 
                           => eshift_19_port);
   C2382 : GTECH_XOR2 port map( A => p_plane_45_port, B => p_plane_36_port, Z 
                           => eshift_18_port);
   C2383 : GTECH_XOR2 port map( A => p_plane_44_port, B => p_plane_35_port, Z 
                           => eshift_17_port);
   C2384 : GTECH_XOR2 port map( A => p_plane_43_port, B => p_plane_34_port, Z 
                           => eshift_16_port);
   C2385 : GTECH_XOR2 port map( A => p_plane_42_port, B => p_plane_33_port, Z 
                           => eshift_15_port);
   C2386 : GTECH_XOR2 port map( A => p_plane_41_port, B => p_plane_32_port, Z 
                           => eshift_14_port);
   C2387 : GTECH_XOR2 port map( A => p_plane_40_port, B => p_plane_63_port, Z 
                           => eshift_13_port);
   C2388 : GTECH_XOR2 port map( A => p_plane_39_port, B => p_plane_62_port, Z 
                           => eshift_12_port);
   C2389 : GTECH_XOR2 port map( A => p_plane_38_port, B => p_plane_61_port, Z 
                           => eshift_11_port);
   C2390 : GTECH_XOR2 port map( A => p_plane_37_port, B => p_plane_60_port, Z 
                           => eshift_10_port);
   C2391 : GTECH_XOR2 port map( A => p_plane_36_port, B => p_plane_59_port, Z 
                           => eshift_9_port);
   C2392 : GTECH_XOR2 port map( A => p_plane_35_port, B => p_plane_58_port, Z 
                           => eshift_8_port);
   C2393 : GTECH_XOR2 port map( A => p_plane_34_port, B => p_plane_57_port, Z 
                           => eshift_7_port);
   C2394 : GTECH_XOR2 port map( A => p_plane_33_port, B => p_plane_56_port, Z 
                           => eshift_6_port);
   C2395 : GTECH_XOR2 port map( A => p_plane_32_port, B => p_plane_55_port, Z 
                           => eshift_5_port);
   C2396 : GTECH_XOR2 port map( A => p_plane_63_port, B => p_plane_54_port, Z 
                           => eshift_4_port);
   C2397 : GTECH_XOR2 port map( A => p_plane_62_port, B => p_plane_53_port, Z 
                           => eshift_3_port);
   C2398 : GTECH_XOR2 port map( A => p_plane_61_port, B => p_plane_52_port, Z 
                           => eshift_2_port);
   C2399 : GTECH_XOR2 port map( A => p_plane_60_port, B => p_plane_51_port, Z 
                           => eshift_1_port);
   C2400 : GTECH_XOR2 port map( A => p_plane_59_port, B => p_plane_50_port, Z 
                           => eshift_0_port);
   C2401 : GTECH_XOR2 port map( A => INPUT(383), B => eshift_127_port, Z => 
                           plane2_2_127_port);
   C2402 : GTECH_XOR2 port map( A => INPUT(382), B => eshift_126_port, Z => 
                           plane2_2_126_port);
   C2403 : GTECH_XOR2 port map( A => INPUT(381), B => eshift_125_port, Z => 
                           plane2_2_125_port);
   C2404 : GTECH_XOR2 port map( A => INPUT(380), B => eshift_124_port, Z => 
                           plane2_2_124_port);
   C2405 : GTECH_XOR2 port map( A => INPUT(379), B => eshift_123_port, Z => 
                           plane2_2_123_port);
   C2406 : GTECH_XOR2 port map( A => INPUT(378), B => eshift_122_port, Z => 
                           plane2_2_122_port);
   C2407 : GTECH_XOR2 port map( A => INPUT(377), B => eshift_121_port, Z => 
                           plane2_2_121_port);
   C2408 : GTECH_XOR2 port map( A => INPUT(376), B => eshift_120_port, Z => 
                           plane2_2_120_port);
   C2409 : GTECH_XOR2 port map( A => INPUT(375), B => eshift_119_port, Z => 
                           plane2_2_119_port);
   C2410 : GTECH_XOR2 port map( A => INPUT(374), B => eshift_118_port, Z => 
                           plane2_2_118_port);
   C2411 : GTECH_XOR2 port map( A => INPUT(373), B => eshift_117_port, Z => 
                           plane2_2_117_port);
   C2412 : GTECH_XOR2 port map( A => INPUT(372), B => eshift_116_port, Z => 
                           plane2_2_116_port);
   C2413 : GTECH_XOR2 port map( A => INPUT(371), B => eshift_115_port, Z => 
                           plane2_2_115_port);
   C2414 : GTECH_XOR2 port map( A => INPUT(370), B => eshift_114_port, Z => 
                           plane2_2_114_port);
   C2415 : GTECH_XOR2 port map( A => INPUT(369), B => eshift_113_port, Z => 
                           plane2_2_113_port);
   C2416 : GTECH_XOR2 port map( A => INPUT(368), B => eshift_112_port, Z => 
                           plane2_2_112_port);
   C2417 : GTECH_XOR2 port map( A => INPUT(367), B => eshift_111_port, Z => 
                           plane2_2_111_port);
   C2418 : GTECH_XOR2 port map( A => INPUT(366), B => eshift_110_port, Z => 
                           plane2_2_110_port);
   C2419 : GTECH_XOR2 port map( A => INPUT(365), B => eshift_109_port, Z => 
                           plane2_2_109_port);
   C2420 : GTECH_XOR2 port map( A => INPUT(364), B => eshift_108_port, Z => 
                           plane2_2_108_port);
   C2421 : GTECH_XOR2 port map( A => INPUT(363), B => eshift_107_port, Z => 
                           plane2_2_107_port);
   C2422 : GTECH_XOR2 port map( A => INPUT(362), B => eshift_106_port, Z => 
                           plane2_2_106_port);
   C2423 : GTECH_XOR2 port map( A => INPUT(361), B => eshift_105_port, Z => 
                           plane2_2_105_port);
   C2424 : GTECH_XOR2 port map( A => INPUT(360), B => eshift_104_port, Z => 
                           plane2_2_104_port);
   C2425 : GTECH_XOR2 port map( A => INPUT(359), B => eshift_103_port, Z => 
                           plane2_2_103_port);
   C2426 : GTECH_XOR2 port map( A => INPUT(358), B => eshift_102_port, Z => 
                           plane2_2_102_port);
   C2427 : GTECH_XOR2 port map( A => INPUT(357), B => eshift_101_port, Z => 
                           plane2_2_101_port);
   C2428 : GTECH_XOR2 port map( A => INPUT(356), B => eshift_100_port, Z => 
                           plane2_2_100_port);
   C2429 : GTECH_XOR2 port map( A => INPUT(355), B => eshift_99_port, Z => 
                           plane2_2_99_port);
   C2430 : GTECH_XOR2 port map( A => INPUT(354), B => eshift_98_port, Z => 
                           plane2_2_98_port);
   C2431 : GTECH_XOR2 port map( A => INPUT(353), B => eshift_97_port, Z => 
                           plane2_2_97_port);
   C2432 : GTECH_XOR2 port map( A => INPUT(352), B => eshift_96_port, Z => 
                           plane2_2_96_port);
   C2433 : GTECH_XOR2 port map( A => INPUT(351), B => eshift_95_port, Z => 
                           plane2_2_95_port);
   C2434 : GTECH_XOR2 port map( A => INPUT(350), B => eshift_94_port, Z => 
                           plane2_2_94_port);
   C2435 : GTECH_XOR2 port map( A => INPUT(349), B => eshift_93_port, Z => 
                           plane2_2_93_port);
   C2436 : GTECH_XOR2 port map( A => INPUT(348), B => eshift_92_port, Z => 
                           plane2_2_92_port);
   C2437 : GTECH_XOR2 port map( A => INPUT(347), B => eshift_91_port, Z => 
                           plane2_2_91_port);
   C2438 : GTECH_XOR2 port map( A => INPUT(346), B => eshift_90_port, Z => 
                           plane2_2_90_port);
   C2439 : GTECH_XOR2 port map( A => INPUT(345), B => eshift_89_port, Z => 
                           plane2_2_89_port);
   C2440 : GTECH_XOR2 port map( A => INPUT(344), B => eshift_88_port, Z => 
                           plane2_2_88_port);
   C2441 : GTECH_XOR2 port map( A => INPUT(343), B => eshift_87_port, Z => 
                           plane2_2_87_port);
   C2442 : GTECH_XOR2 port map( A => INPUT(342), B => eshift_86_port, Z => 
                           plane2_2_86_port);
   C2443 : GTECH_XOR2 port map( A => INPUT(341), B => eshift_85_port, Z => 
                           plane2_2_85_port);
   C2444 : GTECH_XOR2 port map( A => INPUT(340), B => eshift_84_port, Z => 
                           plane2_2_84_port);
   C2445 : GTECH_XOR2 port map( A => INPUT(339), B => eshift_83_port, Z => 
                           plane2_2_83_port);
   C2446 : GTECH_XOR2 port map( A => INPUT(338), B => eshift_82_port, Z => 
                           plane2_2_82_port);
   C2447 : GTECH_XOR2 port map( A => INPUT(337), B => eshift_81_port, Z => 
                           plane2_2_81_port);
   C2448 : GTECH_XOR2 port map( A => INPUT(336), B => eshift_80_port, Z => 
                           plane2_2_80_port);
   C2449 : GTECH_XOR2 port map( A => INPUT(335), B => eshift_79_port, Z => 
                           plane2_2_79_port);
   C2450 : GTECH_XOR2 port map( A => INPUT(334), B => eshift_78_port, Z => 
                           plane2_2_78_port);
   C2451 : GTECH_XOR2 port map( A => INPUT(333), B => eshift_77_port, Z => 
                           plane2_2_77_port);
   C2452 : GTECH_XOR2 port map( A => INPUT(332), B => eshift_76_port, Z => 
                           plane2_2_76_port);
   C2453 : GTECH_XOR2 port map( A => INPUT(331), B => eshift_75_port, Z => 
                           plane2_2_75_port);
   C2454 : GTECH_XOR2 port map( A => INPUT(330), B => eshift_74_port, Z => 
                           plane2_2_74_port);
   C2455 : GTECH_XOR2 port map( A => INPUT(329), B => eshift_73_port, Z => 
                           plane2_2_73_port);
   C2456 : GTECH_XOR2 port map( A => INPUT(328), B => eshift_72_port, Z => 
                           plane2_2_72_port);
   C2457 : GTECH_XOR2 port map( A => INPUT(327), B => eshift_71_port, Z => 
                           plane2_2_71_port);
   C2458 : GTECH_XOR2 port map( A => INPUT(326), B => eshift_70_port, Z => 
                           plane2_2_70_port);
   C2459 : GTECH_XOR2 port map( A => INPUT(325), B => eshift_69_port, Z => 
                           plane2_2_69_port);
   C2460 : GTECH_XOR2 port map( A => INPUT(324), B => eshift_68_port, Z => 
                           plane2_2_68_port);
   C2461 : GTECH_XOR2 port map( A => INPUT(323), B => eshift_67_port, Z => 
                           plane2_2_67_port);
   C2462 : GTECH_XOR2 port map( A => INPUT(322), B => eshift_66_port, Z => 
                           plane2_2_66_port);
   C2463 : GTECH_XOR2 port map( A => INPUT(321), B => eshift_65_port, Z => 
                           plane2_2_65_port);
   C2464 : GTECH_XOR2 port map( A => INPUT(320), B => eshift_64_port, Z => 
                           plane2_2_64_port);
   C2465 : GTECH_XOR2 port map( A => INPUT(319), B => eshift_63_port, Z => 
                           plane2_2_63_port);
   C2466 : GTECH_XOR2 port map( A => INPUT(318), B => eshift_62_port, Z => 
                           plane2_2_62_port);
   C2467 : GTECH_XOR2 port map( A => INPUT(317), B => eshift_61_port, Z => 
                           plane2_2_61_port);
   C2468 : GTECH_XOR2 port map( A => INPUT(316), B => eshift_60_port, Z => 
                           plane2_2_60_port);
   C2469 : GTECH_XOR2 port map( A => INPUT(315), B => eshift_59_port, Z => 
                           plane2_2_59_port);
   C2470 : GTECH_XOR2 port map( A => INPUT(314), B => eshift_58_port, Z => 
                           plane2_2_58_port);
   C2471 : GTECH_XOR2 port map( A => INPUT(313), B => eshift_57_port, Z => 
                           plane2_2_57_port);
   C2472 : GTECH_XOR2 port map( A => INPUT(312), B => eshift_56_port, Z => 
                           plane2_2_56_port);
   C2473 : GTECH_XOR2 port map( A => INPUT(311), B => eshift_55_port, Z => 
                           plane2_2_55_port);
   C2474 : GTECH_XOR2 port map( A => INPUT(310), B => eshift_54_port, Z => 
                           plane2_2_54_port);
   C2475 : GTECH_XOR2 port map( A => INPUT(309), B => eshift_53_port, Z => 
                           plane2_2_53_port);
   C2476 : GTECH_XOR2 port map( A => INPUT(308), B => eshift_52_port, Z => 
                           plane2_2_52_port);
   C2477 : GTECH_XOR2 port map( A => INPUT(307), B => eshift_51_port, Z => 
                           plane2_2_51_port);
   C2478 : GTECH_XOR2 port map( A => INPUT(306), B => eshift_50_port, Z => 
                           plane2_2_50_port);
   C2479 : GTECH_XOR2 port map( A => INPUT(305), B => eshift_49_port, Z => 
                           plane2_2_49_port);
   C2480 : GTECH_XOR2 port map( A => INPUT(304), B => eshift_48_port, Z => 
                           plane2_2_48_port);
   C2481 : GTECH_XOR2 port map( A => INPUT(303), B => eshift_47_port, Z => 
                           plane2_2_47_port);
   C2482 : GTECH_XOR2 port map( A => INPUT(302), B => eshift_46_port, Z => 
                           plane2_2_46_port);
   C2483 : GTECH_XOR2 port map( A => INPUT(301), B => eshift_45_port, Z => 
                           plane2_2_45_port);
   C2484 : GTECH_XOR2 port map( A => INPUT(300), B => eshift_44_port, Z => 
                           plane2_2_44_port);
   C2485 : GTECH_XOR2 port map( A => INPUT(299), B => eshift_43_port, Z => 
                           plane2_2_43_port);
   C2486 : GTECH_XOR2 port map( A => INPUT(298), B => eshift_42_port, Z => 
                           plane2_2_42_port);
   C2487 : GTECH_XOR2 port map( A => INPUT(297), B => eshift_41_port, Z => 
                           plane2_2_41_port);
   C2488 : GTECH_XOR2 port map( A => INPUT(296), B => eshift_40_port, Z => 
                           plane2_2_40_port);
   C2489 : GTECH_XOR2 port map( A => INPUT(295), B => eshift_39_port, Z => 
                           plane2_2_39_port);
   C2490 : GTECH_XOR2 port map( A => INPUT(294), B => eshift_38_port, Z => 
                           plane2_2_38_port);
   C2491 : GTECH_XOR2 port map( A => INPUT(293), B => eshift_37_port, Z => 
                           plane2_2_37_port);
   C2492 : GTECH_XOR2 port map( A => INPUT(292), B => eshift_36_port, Z => 
                           plane2_2_36_port);
   C2493 : GTECH_XOR2 port map( A => INPUT(291), B => eshift_35_port, Z => 
                           plane2_2_35_port);
   C2494 : GTECH_XOR2 port map( A => INPUT(290), B => eshift_34_port, Z => 
                           plane2_2_34_port);
   C2495 : GTECH_XOR2 port map( A => INPUT(289), B => eshift_33_port, Z => 
                           plane2_2_33_port);
   C2496 : GTECH_XOR2 port map( A => INPUT(288), B => eshift_32_port, Z => 
                           plane2_2_32_port);
   C2497 : GTECH_XOR2 port map( A => INPUT(287), B => eshift_31_port, Z => 
                           plane2_2_31_port);
   C2498 : GTECH_XOR2 port map( A => INPUT(286), B => eshift_30_port, Z => 
                           plane2_2_30_port);
   C2499 : GTECH_XOR2 port map( A => INPUT(285), B => eshift_29_port, Z => 
                           plane2_2_29_port);
   C2500 : GTECH_XOR2 port map( A => INPUT(284), B => eshift_28_port, Z => 
                           plane2_2_28_port);
   C2501 : GTECH_XOR2 port map( A => INPUT(283), B => eshift_27_port, Z => 
                           plane2_2_27_port);
   C2502 : GTECH_XOR2 port map( A => INPUT(282), B => eshift_26_port, Z => 
                           plane2_2_26_port);
   C2503 : GTECH_XOR2 port map( A => INPUT(281), B => eshift_25_port, Z => 
                           plane2_2_25_port);
   C2504 : GTECH_XOR2 port map( A => INPUT(280), B => eshift_24_port, Z => 
                           plane2_2_24_port);
   C2505 : GTECH_XOR2 port map( A => INPUT(279), B => eshift_23_port, Z => 
                           plane2_2_23_port);
   C2506 : GTECH_XOR2 port map( A => INPUT(278), B => eshift_22_port, Z => 
                           plane2_2_22_port);
   C2507 : GTECH_XOR2 port map( A => INPUT(277), B => eshift_21_port, Z => 
                           plane2_2_21_port);
   C2508 : GTECH_XOR2 port map( A => INPUT(276), B => eshift_20_port, Z => 
                           plane2_2_20_port);
   C2509 : GTECH_XOR2 port map( A => INPUT(275), B => eshift_19_port, Z => 
                           plane2_2_19_port);
   C2510 : GTECH_XOR2 port map( A => INPUT(274), B => eshift_18_port, Z => 
                           plane2_2_18_port);
   C2511 : GTECH_XOR2 port map( A => INPUT(273), B => eshift_17_port, Z => 
                           plane2_2_17_port);
   C2512 : GTECH_XOR2 port map( A => INPUT(272), B => eshift_16_port, Z => 
                           plane2_2_16_port);
   C2513 : GTECH_XOR2 port map( A => INPUT(271), B => eshift_15_port, Z => 
                           plane2_2_15_port);
   C2514 : GTECH_XOR2 port map( A => INPUT(270), B => eshift_14_port, Z => 
                           plane2_2_14_port);
   C2515 : GTECH_XOR2 port map( A => INPUT(269), B => eshift_13_port, Z => 
                           plane2_2_13_port);
   C2516 : GTECH_XOR2 port map( A => INPUT(268), B => eshift_12_port, Z => 
                           plane2_2_12_port);
   C2517 : GTECH_XOR2 port map( A => INPUT(267), B => eshift_11_port, Z => 
                           plane2_2_11_port);
   C2518 : GTECH_XOR2 port map( A => INPUT(266), B => eshift_10_port, Z => 
                           plane2_2_10_port);
   C2519 : GTECH_XOR2 port map( A => INPUT(265), B => eshift_9_port, Z => 
                           plane2_2_9_port);
   C2520 : GTECH_XOR2 port map( A => INPUT(264), B => eshift_8_port, Z => 
                           plane2_2_8_port);
   C2521 : GTECH_XOR2 port map( A => INPUT(263), B => eshift_7_port, Z => 
                           plane2_2_7_port);
   C2522 : GTECH_XOR2 port map( A => INPUT(262), B => eshift_6_port, Z => 
                           plane2_2_6_port);
   C2523 : GTECH_XOR2 port map( A => INPUT(261), B => eshift_5_port, Z => 
                           plane2_2_5_port);
   C2524 : GTECH_XOR2 port map( A => INPUT(260), B => eshift_4_port, Z => 
                           plane2_2_4_port);
   C2525 : GTECH_XOR2 port map( A => INPUT(259), B => eshift_3_port, Z => 
                           plane2_2_3_port);
   C2526 : GTECH_XOR2 port map( A => INPUT(258), B => eshift_2_port, Z => 
                           plane2_2_2_port);
   C2527 : GTECH_XOR2 port map( A => INPUT(257), B => eshift_1_port, Z => 
                           plane2_2_1_port);
   C2528 : GTECH_XOR2 port map( A => INPUT(256), B => eshift_0_port, Z => 
                           plane2_2_0_port);
   C2529 : GTECH_XOR2 port map( A => INPUT(255), B => eshift_127_port, Z => 
                           plane1_2_127_port);
   C2530 : GTECH_XOR2 port map( A => INPUT(254), B => eshift_126_port, Z => 
                           plane1_2_126_port);
   C2531 : GTECH_XOR2 port map( A => INPUT(253), B => eshift_125_port, Z => 
                           plane1_2_125_port);
   C2532 : GTECH_XOR2 port map( A => INPUT(252), B => eshift_124_port, Z => 
                           plane1_2_124_port);
   C2533 : GTECH_XOR2 port map( A => INPUT(251), B => eshift_123_port, Z => 
                           plane1_2_123_port);
   C2534 : GTECH_XOR2 port map( A => INPUT(250), B => eshift_122_port, Z => 
                           plane1_2_122_port);
   C2535 : GTECH_XOR2 port map( A => INPUT(249), B => eshift_121_port, Z => 
                           plane1_2_121_port);
   C2536 : GTECH_XOR2 port map( A => INPUT(248), B => eshift_120_port, Z => 
                           plane1_2_120_port);
   C2537 : GTECH_XOR2 port map( A => INPUT(247), B => eshift_119_port, Z => 
                           plane1_2_119_port);
   C2538 : GTECH_XOR2 port map( A => INPUT(246), B => eshift_118_port, Z => 
                           plane1_2_118_port);
   C2539 : GTECH_XOR2 port map( A => INPUT(245), B => eshift_117_port, Z => 
                           plane1_2_117_port);
   C2540 : GTECH_XOR2 port map( A => INPUT(244), B => eshift_116_port, Z => 
                           plane1_2_116_port);
   C2541 : GTECH_XOR2 port map( A => INPUT(243), B => eshift_115_port, Z => 
                           plane1_2_115_port);
   C2542 : GTECH_XOR2 port map( A => INPUT(242), B => eshift_114_port, Z => 
                           plane1_2_114_port);
   C2543 : GTECH_XOR2 port map( A => INPUT(241), B => eshift_113_port, Z => 
                           plane1_2_113_port);
   C2544 : GTECH_XOR2 port map( A => INPUT(240), B => eshift_112_port, Z => 
                           plane1_2_112_port);
   C2545 : GTECH_XOR2 port map( A => INPUT(239), B => eshift_111_port, Z => 
                           plane1_2_111_port);
   C2546 : GTECH_XOR2 port map( A => INPUT(238), B => eshift_110_port, Z => 
                           plane1_2_110_port);
   C2547 : GTECH_XOR2 port map( A => INPUT(237), B => eshift_109_port, Z => 
                           plane1_2_109_port);
   C2548 : GTECH_XOR2 port map( A => INPUT(236), B => eshift_108_port, Z => 
                           plane1_2_108_port);
   C2549 : GTECH_XOR2 port map( A => INPUT(235), B => eshift_107_port, Z => 
                           plane1_2_107_port);
   C2550 : GTECH_XOR2 port map( A => INPUT(234), B => eshift_106_port, Z => 
                           plane1_2_106_port);
   C2551 : GTECH_XOR2 port map( A => INPUT(233), B => eshift_105_port, Z => 
                           plane1_2_105_port);
   C2552 : GTECH_XOR2 port map( A => INPUT(232), B => eshift_104_port, Z => 
                           plane1_2_104_port);
   C2553 : GTECH_XOR2 port map( A => INPUT(231), B => eshift_103_port, Z => 
                           plane1_2_103_port);
   C2554 : GTECH_XOR2 port map( A => INPUT(230), B => eshift_102_port, Z => 
                           plane1_2_102_port);
   C2555 : GTECH_XOR2 port map( A => INPUT(229), B => eshift_101_port, Z => 
                           plane1_2_101_port);
   C2556 : GTECH_XOR2 port map( A => INPUT(228), B => eshift_100_port, Z => 
                           plane1_2_100_port);
   C2557 : GTECH_XOR2 port map( A => INPUT(227), B => eshift_99_port, Z => 
                           plane1_2_99_port);
   C2558 : GTECH_XOR2 port map( A => INPUT(226), B => eshift_98_port, Z => 
                           plane1_2_98_port);
   C2559 : GTECH_XOR2 port map( A => INPUT(225), B => eshift_97_port, Z => 
                           plane1_2_97_port);
   C2560 : GTECH_XOR2 port map( A => INPUT(224), B => eshift_96_port, Z => 
                           plane1_2_96_port);
   C2561 : GTECH_XOR2 port map( A => INPUT(223), B => eshift_95_port, Z => 
                           plane1_2_95_port);
   C2562 : GTECH_XOR2 port map( A => INPUT(222), B => eshift_94_port, Z => 
                           plane1_2_94_port);
   C2563 : GTECH_XOR2 port map( A => INPUT(221), B => eshift_93_port, Z => 
                           plane1_2_93_port);
   C2564 : GTECH_XOR2 port map( A => INPUT(220), B => eshift_92_port, Z => 
                           plane1_2_92_port);
   C2565 : GTECH_XOR2 port map( A => INPUT(219), B => eshift_91_port, Z => 
                           plane1_2_91_port);
   C2566 : GTECH_XOR2 port map( A => INPUT(218), B => eshift_90_port, Z => 
                           plane1_2_90_port);
   C2567 : GTECH_XOR2 port map( A => INPUT(217), B => eshift_89_port, Z => 
                           plane1_2_89_port);
   C2568 : GTECH_XOR2 port map( A => INPUT(216), B => eshift_88_port, Z => 
                           plane1_2_88_port);
   C2569 : GTECH_XOR2 port map( A => INPUT(215), B => eshift_87_port, Z => 
                           plane1_2_87_port);
   C2570 : GTECH_XOR2 port map( A => INPUT(214), B => eshift_86_port, Z => 
                           plane1_2_86_port);
   C2571 : GTECH_XOR2 port map( A => INPUT(213), B => eshift_85_port, Z => 
                           plane1_2_85_port);
   C2572 : GTECH_XOR2 port map( A => INPUT(212), B => eshift_84_port, Z => 
                           plane1_2_84_port);
   C2573 : GTECH_XOR2 port map( A => INPUT(211), B => eshift_83_port, Z => 
                           plane1_2_83_port);
   C2574 : GTECH_XOR2 port map( A => INPUT(210), B => eshift_82_port, Z => 
                           plane1_2_82_port);
   C2575 : GTECH_XOR2 port map( A => INPUT(209), B => eshift_81_port, Z => 
                           plane1_2_81_port);
   C2576 : GTECH_XOR2 port map( A => INPUT(208), B => eshift_80_port, Z => 
                           plane1_2_80_port);
   C2577 : GTECH_XOR2 port map( A => INPUT(207), B => eshift_79_port, Z => 
                           plane1_2_79_port);
   C2578 : GTECH_XOR2 port map( A => INPUT(206), B => eshift_78_port, Z => 
                           plane1_2_78_port);
   C2579 : GTECH_XOR2 port map( A => INPUT(205), B => eshift_77_port, Z => 
                           plane1_2_77_port);
   C2580 : GTECH_XOR2 port map( A => INPUT(204), B => eshift_76_port, Z => 
                           plane1_2_76_port);
   C2581 : GTECH_XOR2 port map( A => INPUT(203), B => eshift_75_port, Z => 
                           plane1_2_75_port);
   C2582 : GTECH_XOR2 port map( A => INPUT(202), B => eshift_74_port, Z => 
                           plane1_2_74_port);
   C2583 : GTECH_XOR2 port map( A => INPUT(201), B => eshift_73_port, Z => 
                           plane1_2_73_port);
   C2584 : GTECH_XOR2 port map( A => INPUT(200), B => eshift_72_port, Z => 
                           plane1_2_72_port);
   C2585 : GTECH_XOR2 port map( A => INPUT(199), B => eshift_71_port, Z => 
                           plane1_2_71_port);
   C2586 : GTECH_XOR2 port map( A => INPUT(198), B => eshift_70_port, Z => 
                           plane1_2_70_port);
   C2587 : GTECH_XOR2 port map( A => INPUT(197), B => eshift_69_port, Z => 
                           plane1_2_69_port);
   C2588 : GTECH_XOR2 port map( A => INPUT(196), B => eshift_68_port, Z => 
                           plane1_2_68_port);
   C2589 : GTECH_XOR2 port map( A => INPUT(195), B => eshift_67_port, Z => 
                           plane1_2_67_port);
   C2590 : GTECH_XOR2 port map( A => INPUT(194), B => eshift_66_port, Z => 
                           plane1_2_66_port);
   C2591 : GTECH_XOR2 port map( A => INPUT(193), B => eshift_65_port, Z => 
                           plane1_2_65_port);
   C2592 : GTECH_XOR2 port map( A => INPUT(192), B => eshift_64_port, Z => 
                           plane1_2_64_port);
   C2593 : GTECH_XOR2 port map( A => INPUT(191), B => eshift_63_port, Z => 
                           plane1_2_63_port);
   C2594 : GTECH_XOR2 port map( A => INPUT(190), B => eshift_62_port, Z => 
                           plane1_2_62_port);
   C2595 : GTECH_XOR2 port map( A => INPUT(189), B => eshift_61_port, Z => 
                           plane1_2_61_port);
   C2596 : GTECH_XOR2 port map( A => INPUT(188), B => eshift_60_port, Z => 
                           plane1_2_60_port);
   C2597 : GTECH_XOR2 port map( A => INPUT(187), B => eshift_59_port, Z => 
                           plane1_2_59_port);
   C2598 : GTECH_XOR2 port map( A => INPUT(186), B => eshift_58_port, Z => 
                           plane1_2_58_port);
   C2599 : GTECH_XOR2 port map( A => INPUT(185), B => eshift_57_port, Z => 
                           plane1_2_57_port);
   C2600 : GTECH_XOR2 port map( A => INPUT(184), B => eshift_56_port, Z => 
                           plane1_2_56_port);
   C2601 : GTECH_XOR2 port map( A => INPUT(183), B => eshift_55_port, Z => 
                           plane1_2_55_port);
   C2602 : GTECH_XOR2 port map( A => INPUT(182), B => eshift_54_port, Z => 
                           plane1_2_54_port);
   C2603 : GTECH_XOR2 port map( A => INPUT(181), B => eshift_53_port, Z => 
                           plane1_2_53_port);
   C2604 : GTECH_XOR2 port map( A => INPUT(180), B => eshift_52_port, Z => 
                           plane1_2_52_port);
   C2605 : GTECH_XOR2 port map( A => INPUT(179), B => eshift_51_port, Z => 
                           plane1_2_51_port);
   C2606 : GTECH_XOR2 port map( A => INPUT(178), B => eshift_50_port, Z => 
                           plane1_2_50_port);
   C2607 : GTECH_XOR2 port map( A => INPUT(177), B => eshift_49_port, Z => 
                           plane1_2_49_port);
   C2608 : GTECH_XOR2 port map( A => INPUT(176), B => eshift_48_port, Z => 
                           plane1_2_48_port);
   C2609 : GTECH_XOR2 port map( A => INPUT(175), B => eshift_47_port, Z => 
                           plane1_2_47_port);
   C2610 : GTECH_XOR2 port map( A => INPUT(174), B => eshift_46_port, Z => 
                           plane1_2_46_port);
   C2611 : GTECH_XOR2 port map( A => INPUT(173), B => eshift_45_port, Z => 
                           plane1_2_45_port);
   C2612 : GTECH_XOR2 port map( A => INPUT(172), B => eshift_44_port, Z => 
                           plane1_2_44_port);
   C2613 : GTECH_XOR2 port map( A => INPUT(171), B => eshift_43_port, Z => 
                           plane1_2_43_port);
   C2614 : GTECH_XOR2 port map( A => INPUT(170), B => eshift_42_port, Z => 
                           plane1_2_42_port);
   C2615 : GTECH_XOR2 port map( A => INPUT(169), B => eshift_41_port, Z => 
                           plane1_2_41_port);
   C2616 : GTECH_XOR2 port map( A => INPUT(168), B => eshift_40_port, Z => 
                           plane1_2_40_port);
   C2617 : GTECH_XOR2 port map( A => INPUT(167), B => eshift_39_port, Z => 
                           plane1_2_39_port);
   C2618 : GTECH_XOR2 port map( A => INPUT(166), B => eshift_38_port, Z => 
                           plane1_2_38_port);
   C2619 : GTECH_XOR2 port map( A => INPUT(165), B => eshift_37_port, Z => 
                           plane1_2_37_port);
   C2620 : GTECH_XOR2 port map( A => INPUT(164), B => eshift_36_port, Z => 
                           plane1_2_36_port);
   C2621 : GTECH_XOR2 port map( A => INPUT(163), B => eshift_35_port, Z => 
                           plane1_2_35_port);
   C2622 : GTECH_XOR2 port map( A => INPUT(162), B => eshift_34_port, Z => 
                           plane1_2_34_port);
   C2623 : GTECH_XOR2 port map( A => INPUT(161), B => eshift_33_port, Z => 
                           plane1_2_33_port);
   C2624 : GTECH_XOR2 port map( A => INPUT(160), B => eshift_32_port, Z => 
                           plane1_2_32_port);
   C2625 : GTECH_XOR2 port map( A => INPUT(159), B => eshift_31_port, Z => 
                           plane1_2_31_port);
   C2626 : GTECH_XOR2 port map( A => INPUT(158), B => eshift_30_port, Z => 
                           plane1_2_30_port);
   C2627 : GTECH_XOR2 port map( A => INPUT(157), B => eshift_29_port, Z => 
                           plane1_2_29_port);
   C2628 : GTECH_XOR2 port map( A => INPUT(156), B => eshift_28_port, Z => 
                           plane1_2_28_port);
   C2629 : GTECH_XOR2 port map( A => INPUT(155), B => eshift_27_port, Z => 
                           plane1_2_27_port);
   C2630 : GTECH_XOR2 port map( A => INPUT(154), B => eshift_26_port, Z => 
                           plane1_2_26_port);
   C2631 : GTECH_XOR2 port map( A => INPUT(153), B => eshift_25_port, Z => 
                           plane1_2_25_port);
   C2632 : GTECH_XOR2 port map( A => INPUT(152), B => eshift_24_port, Z => 
                           plane1_2_24_port);
   C2633 : GTECH_XOR2 port map( A => INPUT(151), B => eshift_23_port, Z => 
                           plane1_2_23_port);
   C2634 : GTECH_XOR2 port map( A => INPUT(150), B => eshift_22_port, Z => 
                           plane1_2_22_port);
   C2635 : GTECH_XOR2 port map( A => INPUT(149), B => eshift_21_port, Z => 
                           plane1_2_21_port);
   C2636 : GTECH_XOR2 port map( A => INPUT(148), B => eshift_20_port, Z => 
                           plane1_2_20_port);
   C2637 : GTECH_XOR2 port map( A => INPUT(147), B => eshift_19_port, Z => 
                           plane1_2_19_port);
   C2638 : GTECH_XOR2 port map( A => INPUT(146), B => eshift_18_port, Z => 
                           plane1_2_18_port);
   C2639 : GTECH_XOR2 port map( A => INPUT(145), B => eshift_17_port, Z => 
                           plane1_2_17_port);
   C2640 : GTECH_XOR2 port map( A => INPUT(144), B => eshift_16_port, Z => 
                           plane1_2_16_port);
   C2641 : GTECH_XOR2 port map( A => INPUT(143), B => eshift_15_port, Z => 
                           plane1_2_15_port);
   C2642 : GTECH_XOR2 port map( A => INPUT(142), B => eshift_14_port, Z => 
                           plane1_2_14_port);
   C2643 : GTECH_XOR2 port map( A => INPUT(141), B => eshift_13_port, Z => 
                           plane1_2_13_port);
   C2644 : GTECH_XOR2 port map( A => INPUT(140), B => eshift_12_port, Z => 
                           plane1_2_12_port);
   C2645 : GTECH_XOR2 port map( A => INPUT(139), B => eshift_11_port, Z => 
                           plane1_2_11_port);
   C2646 : GTECH_XOR2 port map( A => INPUT(138), B => eshift_10_port, Z => 
                           plane1_2_10_port);
   C2647 : GTECH_XOR2 port map( A => INPUT(137), B => eshift_9_port, Z => 
                           plane1_2_9_port);
   C2648 : GTECH_XOR2 port map( A => INPUT(136), B => eshift_8_port, Z => 
                           plane1_2_8_port);
   C2649 : GTECH_XOR2 port map( A => INPUT(135), B => eshift_7_port, Z => 
                           plane1_2_7_port);
   C2650 : GTECH_XOR2 port map( A => INPUT(134), B => eshift_6_port, Z => 
                           plane1_2_6_port);
   C2651 : GTECH_XOR2 port map( A => INPUT(133), B => eshift_5_port, Z => 
                           plane1_2_5_port);
   C2652 : GTECH_XOR2 port map( A => INPUT(132), B => eshift_4_port, Z => 
                           plane1_2_4_port);
   C2653 : GTECH_XOR2 port map( A => INPUT(131), B => eshift_3_port, Z => 
                           plane1_2_3_port);
   C2654 : GTECH_XOR2 port map( A => INPUT(130), B => eshift_2_port, Z => 
                           plane1_2_2_port);
   C2655 : GTECH_XOR2 port map( A => INPUT(129), B => eshift_1_port, Z => 
                           plane1_2_1_port);
   C2656 : GTECH_XOR2 port map( A => INPUT(128), B => eshift_0_port, Z => 
                           plane1_2_0_port);
   C2657 : GTECH_XOR2 port map( A => INPUT(127), B => eshift_127_port, Z => 
                           plane0_2_127_port);
   C2658 : GTECH_XOR2 port map( A => INPUT(126), B => eshift_126_port, Z => 
                           plane0_2_126_port);
   C2659 : GTECH_XOR2 port map( A => INPUT(125), B => eshift_125_port, Z => 
                           plane0_2_125_port);
   C2660 : GTECH_XOR2 port map( A => INPUT(124), B => eshift_124_port, Z => 
                           plane0_2_124_port);
   C2661 : GTECH_XOR2 port map( A => INPUT(123), B => eshift_123_port, Z => 
                           plane0_2_123_port);
   C2662 : GTECH_XOR2 port map( A => INPUT(122), B => eshift_122_port, Z => 
                           plane0_2_122_port);
   C2663 : GTECH_XOR2 port map( A => INPUT(121), B => eshift_121_port, Z => 
                           plane0_2_121_port);
   C2664 : GTECH_XOR2 port map( A => INPUT(120), B => eshift_120_port, Z => 
                           plane0_2_120_port);
   C2665 : GTECH_XOR2 port map( A => INPUT(119), B => eshift_119_port, Z => 
                           plane0_2_119_port);
   C2666 : GTECH_XOR2 port map( A => INPUT(118), B => eshift_118_port, Z => 
                           plane0_2_118_port);
   C2667 : GTECH_XOR2 port map( A => INPUT(117), B => eshift_117_port, Z => 
                           plane0_2_117_port);
   C2668 : GTECH_XOR2 port map( A => INPUT(116), B => eshift_116_port, Z => 
                           plane0_2_116_port);
   C2669 : GTECH_XOR2 port map( A => INPUT(115), B => eshift_115_port, Z => 
                           plane0_2_115_port);
   C2670 : GTECH_XOR2 port map( A => INPUT(114), B => eshift_114_port, Z => 
                           plane0_2_114_port);
   C2671 : GTECH_XOR2 port map( A => INPUT(113), B => eshift_113_port, Z => 
                           plane0_2_113_port);
   C2672 : GTECH_XOR2 port map( A => INPUT(112), B => eshift_112_port, Z => 
                           plane0_2_112_port);
   C2673 : GTECH_XOR2 port map( A => INPUT(111), B => eshift_111_port, Z => 
                           plane0_2_111_port);
   C2674 : GTECH_XOR2 port map( A => INPUT(110), B => eshift_110_port, Z => 
                           plane0_2_110_port);
   C2675 : GTECH_XOR2 port map( A => INPUT(109), B => eshift_109_port, Z => 
                           plane0_2_109_port);
   C2676 : GTECH_XOR2 port map( A => INPUT(108), B => eshift_108_port, Z => 
                           plane0_2_108_port);
   C2677 : GTECH_XOR2 port map( A => INPUT(107), B => eshift_107_port, Z => 
                           plane0_2_107_port);
   C2678 : GTECH_XOR2 port map( A => INPUT(106), B => eshift_106_port, Z => 
                           plane0_2_106_port);
   C2679 : GTECH_XOR2 port map( A => INPUT(105), B => eshift_105_port, Z => 
                           plane0_2_105_port);
   C2680 : GTECH_XOR2 port map( A => INPUT(104), B => eshift_104_port, Z => 
                           plane0_2_104_port);
   C2681 : GTECH_XOR2 port map( A => INPUT(103), B => eshift_103_port, Z => 
                           plane0_2_103_port);
   C2682 : GTECH_XOR2 port map( A => INPUT(102), B => eshift_102_port, Z => 
                           plane0_2_102_port);
   C2683 : GTECH_XOR2 port map( A => INPUT(101), B => eshift_101_port, Z => 
                           plane0_2_101_port);
   C2684 : GTECH_XOR2 port map( A => INPUT(100), B => eshift_100_port, Z => 
                           plane0_2_100_port);
   C2685 : GTECH_XOR2 port map( A => INPUT(99), B => eshift_99_port, Z => 
                           plane0_2_99_port);
   C2686 : GTECH_XOR2 port map( A => INPUT(98), B => eshift_98_port, Z => 
                           plane0_2_98_port);
   C2687 : GTECH_XOR2 port map( A => INPUT(97), B => eshift_97_port, Z => 
                           plane0_2_97_port);
   C2688 : GTECH_XOR2 port map( A => INPUT(96), B => eshift_96_port, Z => 
                           plane0_2_96_port);
   C2689 : GTECH_XOR2 port map( A => INPUT(95), B => eshift_95_port, Z => 
                           plane0_2_95_port);
   C2690 : GTECH_XOR2 port map( A => INPUT(94), B => eshift_94_port, Z => 
                           plane0_2_94_port);
   C2691 : GTECH_XOR2 port map( A => INPUT(93), B => eshift_93_port, Z => 
                           plane0_2_93_port);
   C2692 : GTECH_XOR2 port map( A => INPUT(92), B => eshift_92_port, Z => 
                           plane0_2_92_port);
   C2693 : GTECH_XOR2 port map( A => INPUT(91), B => eshift_91_port, Z => 
                           plane0_2_91_port);
   C2694 : GTECH_XOR2 port map( A => INPUT(90), B => eshift_90_port, Z => 
                           plane0_2_90_port);
   C2695 : GTECH_XOR2 port map( A => INPUT(89), B => eshift_89_port, Z => 
                           plane0_2_89_port);
   C2696 : GTECH_XOR2 port map( A => INPUT(88), B => eshift_88_port, Z => 
                           plane0_2_88_port);
   C2697 : GTECH_XOR2 port map( A => INPUT(87), B => eshift_87_port, Z => 
                           plane0_2_87_port);
   C2698 : GTECH_XOR2 port map( A => INPUT(86), B => eshift_86_port, Z => 
                           plane0_2_86_port);
   C2699 : GTECH_XOR2 port map( A => INPUT(85), B => eshift_85_port, Z => 
                           plane0_2_85_port);
   C2700 : GTECH_XOR2 port map( A => INPUT(84), B => eshift_84_port, Z => 
                           plane0_2_84_port);
   C2701 : GTECH_XOR2 port map( A => INPUT(83), B => eshift_83_port, Z => 
                           plane0_2_83_port);
   C2702 : GTECH_XOR2 port map( A => INPUT(82), B => eshift_82_port, Z => 
                           plane0_2_82_port);
   C2703 : GTECH_XOR2 port map( A => INPUT(81), B => eshift_81_port, Z => 
                           plane0_2_81_port);
   C2704 : GTECH_XOR2 port map( A => INPUT(80), B => eshift_80_port, Z => 
                           plane0_2_80_port);
   C2705 : GTECH_XOR2 port map( A => INPUT(79), B => eshift_79_port, Z => 
                           plane0_2_79_port);
   C2706 : GTECH_XOR2 port map( A => INPUT(78), B => eshift_78_port, Z => 
                           plane0_2_78_port);
   C2707 : GTECH_XOR2 port map( A => INPUT(77), B => eshift_77_port, Z => 
                           plane0_2_77_port);
   C2708 : GTECH_XOR2 port map( A => INPUT(76), B => eshift_76_port, Z => 
                           plane0_2_76_port);
   C2709 : GTECH_XOR2 port map( A => INPUT(75), B => eshift_75_port, Z => 
                           plane0_2_75_port);
   C2710 : GTECH_XOR2 port map( A => INPUT(74), B => eshift_74_port, Z => 
                           plane0_2_74_port);
   C2711 : GTECH_XOR2 port map( A => INPUT(73), B => eshift_73_port, Z => 
                           plane0_2_73_port);
   C2712 : GTECH_XOR2 port map( A => INPUT(72), B => eshift_72_port, Z => 
                           plane0_2_72_port);
   C2713 : GTECH_XOR2 port map( A => INPUT(71), B => eshift_71_port, Z => 
                           plane0_2_71_port);
   C2714 : GTECH_XOR2 port map( A => INPUT(70), B => eshift_70_port, Z => 
                           plane0_2_70_port);
   C2715 : GTECH_XOR2 port map( A => INPUT(69), B => eshift_69_port, Z => 
                           plane0_2_69_port);
   C2716 : GTECH_XOR2 port map( A => INPUT(68), B => eshift_68_port, Z => 
                           plane0_2_68_port);
   C2717 : GTECH_XOR2 port map( A => INPUT(67), B => eshift_67_port, Z => 
                           plane0_2_67_port);
   C2718 : GTECH_XOR2 port map( A => INPUT(66), B => eshift_66_port, Z => 
                           plane0_2_66_port);
   C2719 : GTECH_XOR2 port map( A => INPUT(65), B => eshift_65_port, Z => 
                           plane0_2_65_port);
   C2720 : GTECH_XOR2 port map( A => INPUT(64), B => eshift_64_port, Z => 
                           plane0_2_64_port);
   C2721 : GTECH_XOR2 port map( A => INPUT(63), B => eshift_63_port, Z => 
                           plane0_2_63_port);
   C2722 : GTECH_XOR2 port map( A => INPUT(62), B => eshift_62_port, Z => 
                           plane0_2_62_port);
   C2723 : GTECH_XOR2 port map( A => INPUT(61), B => eshift_61_port, Z => 
                           plane0_2_61_port);
   C2724 : GTECH_XOR2 port map( A => INPUT(60), B => eshift_60_port, Z => 
                           plane0_2_60_port);
   C2725 : GTECH_XOR2 port map( A => INPUT(59), B => eshift_59_port, Z => 
                           plane0_2_59_port);
   C2726 : GTECH_XOR2 port map( A => INPUT(58), B => eshift_58_port, Z => 
                           plane0_2_58_port);
   C2727 : GTECH_XOR2 port map( A => INPUT(57), B => eshift_57_port, Z => 
                           plane0_2_57_port);
   C2728 : GTECH_XOR2 port map( A => INPUT(56), B => eshift_56_port, Z => 
                           plane0_2_56_port);
   C2729 : GTECH_XOR2 port map( A => INPUT(55), B => eshift_55_port, Z => 
                           plane0_2_55_port);
   C2730 : GTECH_XOR2 port map( A => INPUT(54), B => eshift_54_port, Z => 
                           plane0_2_54_port);
   C2731 : GTECH_XOR2 port map( A => INPUT(53), B => eshift_53_port, Z => 
                           plane0_2_53_port);
   C2732 : GTECH_XOR2 port map( A => INPUT(52), B => eshift_52_port, Z => 
                           plane0_2_52_port);
   C2733 : GTECH_XOR2 port map( A => INPUT(51), B => eshift_51_port, Z => 
                           plane0_2_51_port);
   C2734 : GTECH_XOR2 port map( A => INPUT(50), B => eshift_50_port, Z => 
                           plane0_2_50_port);
   C2735 : GTECH_XOR2 port map( A => INPUT(49), B => eshift_49_port, Z => 
                           plane0_2_49_port);
   C2736 : GTECH_XOR2 port map( A => INPUT(48), B => eshift_48_port, Z => 
                           plane0_2_48_port);
   C2737 : GTECH_XOR2 port map( A => INPUT(47), B => eshift_47_port, Z => 
                           plane0_2_47_port);
   C2738 : GTECH_XOR2 port map( A => INPUT(46), B => eshift_46_port, Z => 
                           plane0_2_46_port);
   C2739 : GTECH_XOR2 port map( A => INPUT(45), B => eshift_45_port, Z => 
                           plane0_2_45_port);
   C2740 : GTECH_XOR2 port map( A => INPUT(44), B => eshift_44_port, Z => 
                           plane0_2_44_port);
   C2741 : GTECH_XOR2 port map( A => INPUT(43), B => eshift_43_port, Z => 
                           plane0_2_43_port);
   C2742 : GTECH_XOR2 port map( A => INPUT(42), B => eshift_42_port, Z => 
                           plane0_2_42_port);
   C2743 : GTECH_XOR2 port map( A => INPUT(41), B => eshift_41_port, Z => 
                           plane0_2_41_port);
   C2744 : GTECH_XOR2 port map( A => INPUT(40), B => eshift_40_port, Z => 
                           plane0_2_40_port);
   C2745 : GTECH_XOR2 port map( A => INPUT(39), B => eshift_39_port, Z => 
                           plane0_2_39_port);
   C2746 : GTECH_XOR2 port map( A => INPUT(38), B => eshift_38_port, Z => 
                           plane0_2_38_port);
   C2747 : GTECH_XOR2 port map( A => INPUT(37), B => eshift_37_port, Z => 
                           plane0_2_37_port);
   C2748 : GTECH_XOR2 port map( A => INPUT(36), B => eshift_36_port, Z => 
                           plane0_2_36_port);
   C2749 : GTECH_XOR2 port map( A => INPUT(35), B => eshift_35_port, Z => 
                           plane0_2_35_port);
   C2750 : GTECH_XOR2 port map( A => INPUT(34), B => eshift_34_port, Z => 
                           plane0_2_34_port);
   C2751 : GTECH_XOR2 port map( A => INPUT(33), B => eshift_33_port, Z => 
                           plane0_2_33_port);
   C2752 : GTECH_XOR2 port map( A => INPUT(32), B => eshift_32_port, Z => 
                           plane0_2_32_port);
   C2753 : GTECH_XOR2 port map( A => INPUT(31), B => eshift_31_port, Z => 
                           plane0_2_31_port);
   C2754 : GTECH_XOR2 port map( A => INPUT(30), B => eshift_30_port, Z => 
                           plane0_2_30_port);
   C2755 : GTECH_XOR2 port map( A => INPUT(29), B => eshift_29_port, Z => 
                           plane0_2_29_port);
   C2756 : GTECH_XOR2 port map( A => INPUT(28), B => eshift_28_port, Z => 
                           plane0_2_28_port);
   C2757 : GTECH_XOR2 port map( A => INPUT(27), B => eshift_27_port, Z => 
                           plane0_2_27_port);
   C2758 : GTECH_XOR2 port map( A => INPUT(26), B => eshift_26_port, Z => 
                           plane0_2_26_port);
   C2759 : GTECH_XOR2 port map( A => INPUT(25), B => eshift_25_port, Z => 
                           plane0_2_25_port);
   C2760 : GTECH_XOR2 port map( A => INPUT(24), B => eshift_24_port, Z => 
                           plane0_2_24_port);
   C2761 : GTECH_XOR2 port map( A => INPUT(23), B => eshift_23_port, Z => 
                           plane0_2_23_port);
   C2762 : GTECH_XOR2 port map( A => INPUT(22), B => eshift_22_port, Z => 
                           plane0_2_22_port);
   C2763 : GTECH_XOR2 port map( A => INPUT(21), B => eshift_21_port, Z => 
                           plane0_2_21_port);
   C2764 : GTECH_XOR2 port map( A => INPUT(20), B => eshift_20_port, Z => 
                           plane0_2_20_port);
   C2765 : GTECH_XOR2 port map( A => INPUT(19), B => eshift_19_port, Z => 
                           plane0_2_19_port);
   C2766 : GTECH_XOR2 port map( A => INPUT(18), B => eshift_18_port, Z => 
                           plane0_2_18_port);
   C2767 : GTECH_XOR2 port map( A => INPUT(17), B => eshift_17_port, Z => 
                           plane0_2_17_port);
   C2768 : GTECH_XOR2 port map( A => INPUT(16), B => eshift_16_port, Z => 
                           plane0_2_16_port);
   C2769 : GTECH_XOR2 port map( A => INPUT(15), B => eshift_15_port, Z => 
                           plane0_2_15_port);
   C2770 : GTECH_XOR2 port map( A => INPUT(14), B => eshift_14_port, Z => 
                           plane0_2_14_port);
   C2771 : GTECH_XOR2 port map( A => INPUT(13), B => eshift_13_port, Z => 
                           plane0_2_13_port);
   C2772 : GTECH_XOR2 port map( A => INPUT(12), B => eshift_12_port, Z => 
                           plane0_2_12_port);
   C2773 : GTECH_XOR2 port map( A => INPUT(11), B => eshift_11_port, Z => 
                           plane0_2_11_port);
   C2774 : GTECH_XOR2 port map( A => INPUT(10), B => eshift_10_port, Z => 
                           plane0_2_10_port);
   C2775 : GTECH_XOR2 port map( A => INPUT(9), B => eshift_9_port, Z => 
                           plane0_2_9_port);
   C2776 : GTECH_XOR2 port map( A => INPUT(8), B => eshift_8_port, Z => 
                           plane0_2_8_port);
   C2777 : GTECH_XOR2 port map( A => INPUT(7), B => eshift_7_port, Z => 
                           plane0_2_7_port);
   C2778 : GTECH_XOR2 port map( A => INPUT(6), B => eshift_6_port, Z => 
                           plane0_2_6_port);
   C2779 : GTECH_XOR2 port map( A => INPUT(5), B => eshift_5_port, Z => 
                           plane0_2_5_port);
   C2780 : GTECH_XOR2 port map( A => INPUT(4), B => eshift_4_port, Z => 
                           plane0_2_4_port);
   C2781 : GTECH_XOR2 port map( A => INPUT(3), B => eshift_3_port, Z => 
                           plane0_2_3_port);
   C2782 : GTECH_XOR2 port map( A => INPUT(2), B => eshift_2_port, Z => 
                           plane0_2_2_port);
   C2783 : GTECH_XOR2 port map( A => INPUT(1), B => eshift_1_port, Z => 
                           plane0_2_1_port);
   C2784 : GTECH_XOR2 port map( A => INPUT(0), B => eshift_0_port, Z => 
                           plane0_2_0_port);
   C2785 : GTECH_XOR2 port map( A => plane0_2_107_port, B => X_Logic0_port, Z 
                           => add_rnd_const_small_11_port);
   C2786 : GTECH_XOR2 port map( A => plane0_2_106_port, B => X_Logic0_port, Z 
                           => add_rnd_const_small_10_port);
   C2787 : GTECH_XOR2 port map( A => plane0_2_105_port, B => N172, Z => 
                           add_rnd_const_small_9_port);
   C2788 : GTECH_XOR2 port map( A => plane0_2_104_port, B => N173, Z => 
                           add_rnd_const_small_8_port);
   C2789 : GTECH_XOR2 port map( A => plane0_2_103_port, B => N174, Z => 
                           add_rnd_const_small_7_port);
   C2790 : GTECH_XOR2 port map( A => plane0_2_102_port, B => N175, Z => 
                           add_rnd_const_small_6_port);
   C2791 : GTECH_XOR2 port map( A => plane0_2_101_port, B => N176, Z => 
                           add_rnd_const_small_5_port);
   C2792 : GTECH_XOR2 port map( A => plane0_2_100_port, B => N177, Z => 
                           add_rnd_const_small_4_port);
   C2793 : GTECH_XOR2 port map( A => plane0_2_99_port, B => N178, Z => 
                           add_rnd_const_small_3_port);
   C2794 : GTECH_XOR2 port map( A => plane0_2_98_port, B => N179, Z => 
                           add_rnd_const_small_2_port);
   C2795 : GTECH_XOR2 port map( A => plane0_2_97_port, B => N180, Z => 
                           add_rnd_const_small_1_port);
   C2796 : GTECH_XOR2 port map( A => plane0_2_96_port, B => X_Logic0_port, Z =>
                           add_rnd_const_small_0_port);
   I_20 : GTECH_NOT port map( A => plane1_2_31_port, Z => N181);
   I_21 : GTECH_NOT port map( A => plane1_2_30_port, Z => N182);
   I_22 : GTECH_NOT port map( A => plane1_2_29_port, Z => N183);
   I_23 : GTECH_NOT port map( A => plane1_2_28_port, Z => N184);
   I_24 : GTECH_NOT port map( A => plane1_2_27_port, Z => N185);
   I_25 : GTECH_NOT port map( A => plane1_2_26_port, Z => N186);
   I_26 : GTECH_NOT port map( A => plane1_2_25_port, Z => N187);
   I_27 : GTECH_NOT port map( A => plane1_2_24_port, Z => N188);
   I_28 : GTECH_NOT port map( A => plane1_2_23_port, Z => N189);
   I_29 : GTECH_NOT port map( A => plane1_2_22_port, Z => N190);
   I_30 : GTECH_NOT port map( A => plane1_2_21_port, Z => N191);
   I_31 : GTECH_NOT port map( A => plane1_2_20_port, Z => N192);
   I_32 : GTECH_NOT port map( A => plane1_2_19_port, Z => N193);
   I_33 : GTECH_NOT port map( A => plane1_2_18_port, Z => N194);
   I_34 : GTECH_NOT port map( A => plane1_2_17_port, Z => N195);
   I_35 : GTECH_NOT port map( A => plane1_2_16_port, Z => N196);
   I_36 : GTECH_NOT port map( A => plane1_2_15_port, Z => N197);
   I_37 : GTECH_NOT port map( A => plane1_2_14_port, Z => N198);
   I_38 : GTECH_NOT port map( A => plane1_2_13_port, Z => N199);
   I_39 : GTECH_NOT port map( A => plane1_2_12_port, Z => N200);
   I_40 : GTECH_NOT port map( A => plane1_2_11_port, Z => N201);
   I_41 : GTECH_NOT port map( A => plane1_2_10_port, Z => N202);
   I_42 : GTECH_NOT port map( A => plane1_2_9_port, Z => N203);
   I_43 : GTECH_NOT port map( A => plane1_2_8_port, Z => N204);
   I_44 : GTECH_NOT port map( A => plane1_2_7_port, Z => N205);
   I_45 : GTECH_NOT port map( A => plane1_2_6_port, Z => N206);
   I_46 : GTECH_NOT port map( A => plane1_2_5_port, Z => N207);
   I_47 : GTECH_NOT port map( A => plane1_2_4_port, Z => N208);
   I_48 : GTECH_NOT port map( A => plane1_2_3_port, Z => N209);
   I_49 : GTECH_NOT port map( A => plane1_2_2_port, Z => N210);
   I_50 : GTECH_NOT port map( A => plane1_2_1_port, Z => N211);
   I_51 : GTECH_NOT port map( A => plane1_2_0_port, Z => N212);
   I_52 : GTECH_NOT port map( A => plane1_2_127_port, Z => N213);
   I_53 : GTECH_NOT port map( A => plane1_2_126_port, Z => N214);
   I_54 : GTECH_NOT port map( A => plane1_2_125_port, Z => N215);
   I_55 : GTECH_NOT port map( A => plane1_2_124_port, Z => N216);
   I_56 : GTECH_NOT port map( A => plane1_2_123_port, Z => N217);
   I_57 : GTECH_NOT port map( A => plane1_2_122_port, Z => N218);
   I_58 : GTECH_NOT port map( A => plane1_2_121_port, Z => N219);
   I_59 : GTECH_NOT port map( A => plane1_2_120_port, Z => N220);
   I_60 : GTECH_NOT port map( A => plane1_2_119_port, Z => N221);
   I_61 : GTECH_NOT port map( A => plane1_2_118_port, Z => N222);
   I_62 : GTECH_NOT port map( A => plane1_2_117_port, Z => N223);
   I_63 : GTECH_NOT port map( A => plane1_2_116_port, Z => N224);
   I_64 : GTECH_NOT port map( A => plane1_2_115_port, Z => N225);
   I_65 : GTECH_NOT port map( A => plane1_2_114_port, Z => N226);
   I_66 : GTECH_NOT port map( A => plane1_2_113_port, Z => N227);
   I_67 : GTECH_NOT port map( A => plane1_2_112_port, Z => N228);
   I_68 : GTECH_NOT port map( A => plane1_2_111_port, Z => N229);
   I_69 : GTECH_NOT port map( A => plane1_2_110_port, Z => N230);
   I_70 : GTECH_NOT port map( A => plane1_2_109_port, Z => N231);
   I_71 : GTECH_NOT port map( A => plane1_2_108_port, Z => N232);
   I_72 : GTECH_NOT port map( A => plane1_2_107_port, Z => N233);
   I_73 : GTECH_NOT port map( A => plane1_2_106_port, Z => N234);
   I_74 : GTECH_NOT port map( A => plane1_2_105_port, Z => N235);
   I_75 : GTECH_NOT port map( A => plane1_2_104_port, Z => N236);
   I_76 : GTECH_NOT port map( A => plane1_2_103_port, Z => N237);
   I_77 : GTECH_NOT port map( A => plane1_2_102_port, Z => N238);
   I_78 : GTECH_NOT port map( A => plane1_2_101_port, Z => N239);
   I_79 : GTECH_NOT port map( A => plane1_2_100_port, Z => N240);
   I_80 : GTECH_NOT port map( A => plane1_2_99_port, Z => N241);
   I_81 : GTECH_NOT port map( A => plane1_2_98_port, Z => N242);
   I_82 : GTECH_NOT port map( A => plane1_2_97_port, Z => N243);
   I_83 : GTECH_NOT port map( A => plane1_2_96_port, Z => N244);
   I_84 : GTECH_NOT port map( A => plane1_2_95_port, Z => N245);
   I_85 : GTECH_NOT port map( A => plane1_2_94_port, Z => N246);
   I_86 : GTECH_NOT port map( A => plane1_2_93_port, Z => N247);
   I_87 : GTECH_NOT port map( A => plane1_2_92_port, Z => N248);
   I_88 : GTECH_NOT port map( A => plane1_2_91_port, Z => N249);
   I_89 : GTECH_NOT port map( A => plane1_2_90_port, Z => N250);
   I_90 : GTECH_NOT port map( A => plane1_2_89_port, Z => N251);
   I_91 : GTECH_NOT port map( A => plane1_2_88_port, Z => N252);
   I_92 : GTECH_NOT port map( A => plane1_2_87_port, Z => N253);
   I_93 : GTECH_NOT port map( A => plane1_2_86_port, Z => N254);
   I_94 : GTECH_NOT port map( A => plane1_2_85_port, Z => N255);
   I_95 : GTECH_NOT port map( A => plane1_2_84_port, Z => N256);
   I_96 : GTECH_NOT port map( A => plane1_2_83_port, Z => N257);
   I_97 : GTECH_NOT port map( A => plane1_2_82_port, Z => N258);
   I_98 : GTECH_NOT port map( A => plane1_2_81_port, Z => N259);
   I_99 : GTECH_NOT port map( A => plane1_2_80_port, Z => N260);
   I_100 : GTECH_NOT port map( A => plane1_2_79_port, Z => N261);
   I_101 : GTECH_NOT port map( A => plane1_2_78_port, Z => N262);
   I_102 : GTECH_NOT port map( A => plane1_2_77_port, Z => N263);
   I_103 : GTECH_NOT port map( A => plane1_2_76_port, Z => N264);
   I_104 : GTECH_NOT port map( A => plane1_2_75_port, Z => N265);
   I_105 : GTECH_NOT port map( A => plane1_2_74_port, Z => N266);
   I_106 : GTECH_NOT port map( A => plane1_2_73_port, Z => N267);
   I_107 : GTECH_NOT port map( A => plane1_2_72_port, Z => N268);
   I_108 : GTECH_NOT port map( A => plane1_2_71_port, Z => N269);
   I_109 : GTECH_NOT port map( A => plane1_2_70_port, Z => N270);
   I_110 : GTECH_NOT port map( A => plane1_2_69_port, Z => N271);
   I_111 : GTECH_NOT port map( A => plane1_2_68_port, Z => N272);
   I_112 : GTECH_NOT port map( A => plane1_2_67_port, Z => N273);
   I_113 : GTECH_NOT port map( A => plane1_2_66_port, Z => N274);
   I_114 : GTECH_NOT port map( A => plane1_2_65_port, Z => N275);
   I_115 : GTECH_NOT port map( A => plane1_2_64_port, Z => N276);
   I_116 : GTECH_NOT port map( A => plane1_2_63_port, Z => N277);
   I_117 : GTECH_NOT port map( A => plane1_2_62_port, Z => N278);
   I_118 : GTECH_NOT port map( A => plane1_2_61_port, Z => N279);
   I_119 : GTECH_NOT port map( A => plane1_2_60_port, Z => N280);
   I_120 : GTECH_NOT port map( A => plane1_2_59_port, Z => N281);
   I_121 : GTECH_NOT port map( A => plane1_2_58_port, Z => N282);
   I_122 : GTECH_NOT port map( A => plane1_2_57_port, Z => N283);
   I_123 : GTECH_NOT port map( A => plane1_2_56_port, Z => N284);
   I_124 : GTECH_NOT port map( A => plane1_2_55_port, Z => N285);
   I_125 : GTECH_NOT port map( A => plane1_2_54_port, Z => N286);
   I_126 : GTECH_NOT port map( A => plane1_2_53_port, Z => N287);
   I_127 : GTECH_NOT port map( A => plane1_2_52_port, Z => N288);
   I_128 : GTECH_NOT port map( A => plane1_2_51_port, Z => N289);
   I_129 : GTECH_NOT port map( A => plane1_2_50_port, Z => N290);
   I_130 : GTECH_NOT port map( A => plane1_2_49_port, Z => N291);
   I_131 : GTECH_NOT port map( A => plane1_2_48_port, Z => N292);
   I_132 : GTECH_NOT port map( A => plane1_2_47_port, Z => N293);
   I_133 : GTECH_NOT port map( A => plane1_2_46_port, Z => N294);
   I_134 : GTECH_NOT port map( A => plane1_2_45_port, Z => N295);
   I_135 : GTECH_NOT port map( A => plane1_2_44_port, Z => N296);
   I_136 : GTECH_NOT port map( A => plane1_2_43_port, Z => N297);
   I_137 : GTECH_NOT port map( A => plane1_2_42_port, Z => N298);
   I_138 : GTECH_NOT port map( A => plane1_2_41_port, Z => N299);
   I_139 : GTECH_NOT port map( A => plane1_2_40_port, Z => N300);
   I_140 : GTECH_NOT port map( A => plane1_2_39_port, Z => N301);
   I_141 : GTECH_NOT port map( A => plane1_2_38_port, Z => N302);
   I_142 : GTECH_NOT port map( A => plane1_2_37_port, Z => N303);
   I_143 : GTECH_NOT port map( A => plane1_2_36_port, Z => N304);
   I_144 : GTECH_NOT port map( A => plane1_2_35_port, Z => N305);
   I_145 : GTECH_NOT port map( A => plane1_2_34_port, Z => N306);
   I_146 : GTECH_NOT port map( A => plane1_2_33_port, Z => N307);
   I_147 : GTECH_NOT port map( A => plane1_2_32_port, Z => N308);
   C2925 : GTECH_AND2 port map( A => N181, B => plane2_2_116_port, Z => N309);
   C2926 : GTECH_AND2 port map( A => N182, B => plane2_2_115_port, Z => N310);
   C2927 : GTECH_AND2 port map( A => N183, B => plane2_2_114_port, Z => N311);
   C2928 : GTECH_AND2 port map( A => N184, B => plane2_2_113_port, Z => N312);
   C2929 : GTECH_AND2 port map( A => N185, B => plane2_2_112_port, Z => N313);
   C2930 : GTECH_AND2 port map( A => N186, B => plane2_2_111_port, Z => N314);
   C2931 : GTECH_AND2 port map( A => N187, B => plane2_2_110_port, Z => N315);
   C2932 : GTECH_AND2 port map( A => N188, B => plane2_2_109_port, Z => N316);
   C2933 : GTECH_AND2 port map( A => N189, B => plane2_2_108_port, Z => N317);
   C2934 : GTECH_AND2 port map( A => N190, B => plane2_2_107_port, Z => N318);
   C2935 : GTECH_AND2 port map( A => N191, B => plane2_2_106_port, Z => N319);
   C2936 : GTECH_AND2 port map( A => N192, B => plane2_2_105_port, Z => N320);
   C2937 : GTECH_AND2 port map( A => N193, B => plane2_2_104_port, Z => N321);
   C2938 : GTECH_AND2 port map( A => N194, B => plane2_2_103_port, Z => N322);
   C2939 : GTECH_AND2 port map( A => N195, B => plane2_2_102_port, Z => N323);
   C2940 : GTECH_AND2 port map( A => N196, B => plane2_2_101_port, Z => N324);
   C2941 : GTECH_AND2 port map( A => N197, B => plane2_2_100_port, Z => N325);
   C2942 : GTECH_AND2 port map( A => N198, B => plane2_2_99_port, Z => N326);
   C2943 : GTECH_AND2 port map( A => N199, B => plane2_2_98_port, Z => N327);
   C2944 : GTECH_AND2 port map( A => N200, B => plane2_2_97_port, Z => N328);
   C2945 : GTECH_AND2 port map( A => N201, B => plane2_2_96_port, Z => N329);
   C2946 : GTECH_AND2 port map( A => N202, B => plane2_2_127_port, Z => N330);
   C2947 : GTECH_AND2 port map( A => N203, B => plane2_2_126_port, Z => N331);
   C2948 : GTECH_AND2 port map( A => N204, B => plane2_2_125_port, Z => N332);
   C2949 : GTECH_AND2 port map( A => N205, B => plane2_2_124_port, Z => N333);
   C2950 : GTECH_AND2 port map( A => N206, B => plane2_2_123_port, Z => N334);
   C2951 : GTECH_AND2 port map( A => N207, B => plane2_2_122_port, Z => N335);
   C2952 : GTECH_AND2 port map( A => N208, B => plane2_2_121_port, Z => N336);
   C2953 : GTECH_AND2 port map( A => N209, B => plane2_2_120_port, Z => N337);
   C2954 : GTECH_AND2 port map( A => N210, B => plane2_2_119_port, Z => N338);
   C2955 : GTECH_AND2 port map( A => N211, B => plane2_2_118_port, Z => N339);
   C2956 : GTECH_AND2 port map( A => N212, B => plane2_2_117_port, Z => N340);
   C2957 : GTECH_AND2 port map( A => N213, B => plane2_2_84_port, Z => N341);
   C2958 : GTECH_AND2 port map( A => N214, B => plane2_2_83_port, Z => N342);
   C2959 : GTECH_AND2 port map( A => N215, B => plane2_2_82_port, Z => N343);
   C2960 : GTECH_AND2 port map( A => N216, B => plane2_2_81_port, Z => N344);
   C2961 : GTECH_AND2 port map( A => N217, B => plane2_2_80_port, Z => N345);
   C2962 : GTECH_AND2 port map( A => N218, B => plane2_2_79_port, Z => N346);
   C2963 : GTECH_AND2 port map( A => N219, B => plane2_2_78_port, Z => N347);
   C2964 : GTECH_AND2 port map( A => N220, B => plane2_2_77_port, Z => N348);
   C2965 : GTECH_AND2 port map( A => N221, B => plane2_2_76_port, Z => N349);
   C2966 : GTECH_AND2 port map( A => N222, B => plane2_2_75_port, Z => N350);
   C2967 : GTECH_AND2 port map( A => N223, B => plane2_2_74_port, Z => N351);
   C2968 : GTECH_AND2 port map( A => N224, B => plane2_2_73_port, Z => N352);
   C2969 : GTECH_AND2 port map( A => N225, B => plane2_2_72_port, Z => N353);
   C2970 : GTECH_AND2 port map( A => N226, B => plane2_2_71_port, Z => N354);
   C2971 : GTECH_AND2 port map( A => N227, B => plane2_2_70_port, Z => N355);
   C2972 : GTECH_AND2 port map( A => N228, B => plane2_2_69_port, Z => N356);
   C2973 : GTECH_AND2 port map( A => N229, B => plane2_2_68_port, Z => N357);
   C2974 : GTECH_AND2 port map( A => N230, B => plane2_2_67_port, Z => N358);
   C2975 : GTECH_AND2 port map( A => N231, B => plane2_2_66_port, Z => N359);
   C2976 : GTECH_AND2 port map( A => N232, B => plane2_2_65_port, Z => N360);
   C2977 : GTECH_AND2 port map( A => N233, B => plane2_2_64_port, Z => N361);
   C2978 : GTECH_AND2 port map( A => N234, B => plane2_2_95_port, Z => N362);
   C2979 : GTECH_AND2 port map( A => N235, B => plane2_2_94_port, Z => N363);
   C2980 : GTECH_AND2 port map( A => N236, B => plane2_2_93_port, Z => N364);
   C2981 : GTECH_AND2 port map( A => N237, B => plane2_2_92_port, Z => N365);
   C2982 : GTECH_AND2 port map( A => N238, B => plane2_2_91_port, Z => N366);
   C2983 : GTECH_AND2 port map( A => N239, B => plane2_2_90_port, Z => N367);
   C2984 : GTECH_AND2 port map( A => N240, B => plane2_2_89_port, Z => N368);
   C2985 : GTECH_AND2 port map( A => N241, B => plane2_2_88_port, Z => N369);
   C2986 : GTECH_AND2 port map( A => N242, B => plane2_2_87_port, Z => N370);
   C2987 : GTECH_AND2 port map( A => N243, B => plane2_2_86_port, Z => N371);
   C2988 : GTECH_AND2 port map( A => N244, B => plane2_2_85_port, Z => N372);
   C2989 : GTECH_AND2 port map( A => N245, B => plane2_2_52_port, Z => N373);
   C2990 : GTECH_AND2 port map( A => N246, B => plane2_2_51_port, Z => N374);
   C2991 : GTECH_AND2 port map( A => N247, B => plane2_2_50_port, Z => N375);
   C2992 : GTECH_AND2 port map( A => N248, B => plane2_2_49_port, Z => N376);
   C2993 : GTECH_AND2 port map( A => N249, B => plane2_2_48_port, Z => N377);
   C2994 : GTECH_AND2 port map( A => N250, B => plane2_2_47_port, Z => N378);
   C2995 : GTECH_AND2 port map( A => N251, B => plane2_2_46_port, Z => N379);
   C2996 : GTECH_AND2 port map( A => N252, B => plane2_2_45_port, Z => N380);
   C2997 : GTECH_AND2 port map( A => N253, B => plane2_2_44_port, Z => N381);
   C2998 : GTECH_AND2 port map( A => N254, B => plane2_2_43_port, Z => N382);
   C2999 : GTECH_AND2 port map( A => N255, B => plane2_2_42_port, Z => N383);
   C3000 : GTECH_AND2 port map( A => N256, B => plane2_2_41_port, Z => N384);
   C3001 : GTECH_AND2 port map( A => N257, B => plane2_2_40_port, Z => N385);
   C3002 : GTECH_AND2 port map( A => N258, B => plane2_2_39_port, Z => N386);
   C3003 : GTECH_AND2 port map( A => N259, B => plane2_2_38_port, Z => N387);
   C3004 : GTECH_AND2 port map( A => N260, B => plane2_2_37_port, Z => N388);
   C3005 : GTECH_AND2 port map( A => N261, B => plane2_2_36_port, Z => N389);
   C3006 : GTECH_AND2 port map( A => N262, B => plane2_2_35_port, Z => N390);
   C3007 : GTECH_AND2 port map( A => N263, B => plane2_2_34_port, Z => N391);
   C3008 : GTECH_AND2 port map( A => N264, B => plane2_2_33_port, Z => N392);
   C3009 : GTECH_AND2 port map( A => N265, B => plane2_2_32_port, Z => N393);
   C3010 : GTECH_AND2 port map( A => N266, B => plane2_2_63_port, Z => N394);
   C3011 : GTECH_AND2 port map( A => N267, B => plane2_2_62_port, Z => N395);
   C3012 : GTECH_AND2 port map( A => N268, B => plane2_2_61_port, Z => N396);
   C3013 : GTECH_AND2 port map( A => N269, B => plane2_2_60_port, Z => N397);
   C3014 : GTECH_AND2 port map( A => N270, B => plane2_2_59_port, Z => N398);
   C3015 : GTECH_AND2 port map( A => N271, B => plane2_2_58_port, Z => N399);
   C3016 : GTECH_AND2 port map( A => N272, B => plane2_2_57_port, Z => N400);
   C3017 : GTECH_AND2 port map( A => N273, B => plane2_2_56_port, Z => N401);
   C3018 : GTECH_AND2 port map( A => N274, B => plane2_2_55_port, Z => N402);
   C3019 : GTECH_AND2 port map( A => N275, B => plane2_2_54_port, Z => N403);
   C3020 : GTECH_AND2 port map( A => N276, B => plane2_2_53_port, Z => N404);
   C3021 : GTECH_AND2 port map( A => N277, B => plane2_2_20_port, Z => N405);
   C3022 : GTECH_AND2 port map( A => N278, B => plane2_2_19_port, Z => N406);
   C3023 : GTECH_AND2 port map( A => N279, B => plane2_2_18_port, Z => N407);
   C3024 : GTECH_AND2 port map( A => N280, B => plane2_2_17_port, Z => N408);
   C3025 : GTECH_AND2 port map( A => N281, B => plane2_2_16_port, Z => N409);
   C3026 : GTECH_AND2 port map( A => N282, B => plane2_2_15_port, Z => N410);
   C3027 : GTECH_AND2 port map( A => N283, B => plane2_2_14_port, Z => N411);
   C3028 : GTECH_AND2 port map( A => N284, B => plane2_2_13_port, Z => N412);
   C3029 : GTECH_AND2 port map( A => N285, B => plane2_2_12_port, Z => N413);
   C3030 : GTECH_AND2 port map( A => N286, B => plane2_2_11_port, Z => N414);
   C3031 : GTECH_AND2 port map( A => N287, B => plane2_2_10_port, Z => N415);
   C3032 : GTECH_AND2 port map( A => N288, B => plane2_2_9_port, Z => N416);
   C3033 : GTECH_AND2 port map( A => N289, B => plane2_2_8_port, Z => N417);
   C3034 : GTECH_AND2 port map( A => N290, B => plane2_2_7_port, Z => N418);
   C3035 : GTECH_AND2 port map( A => N291, B => plane2_2_6_port, Z => N419);
   C3036 : GTECH_AND2 port map( A => N292, B => plane2_2_5_port, Z => N420);
   C3037 : GTECH_AND2 port map( A => N293, B => plane2_2_4_port, Z => N421);
   C3038 : GTECH_AND2 port map( A => N294, B => plane2_2_3_port, Z => N422);
   C3039 : GTECH_AND2 port map( A => N295, B => plane2_2_2_port, Z => N423);
   C3040 : GTECH_AND2 port map( A => N296, B => plane2_2_1_port, Z => N424);
   C3041 : GTECH_AND2 port map( A => N297, B => plane2_2_0_port, Z => N425);
   C3042 : GTECH_AND2 port map( A => N298, B => plane2_2_31_port, Z => N426);
   C3043 : GTECH_AND2 port map( A => N299, B => plane2_2_30_port, Z => N427);
   C3044 : GTECH_AND2 port map( A => N300, B => plane2_2_29_port, Z => N428);
   C3045 : GTECH_AND2 port map( A => N301, B => plane2_2_28_port, Z => N429);
   C3046 : GTECH_AND2 port map( A => N302, B => plane2_2_27_port, Z => N430);
   C3047 : GTECH_AND2 port map( A => N303, B => plane2_2_26_port, Z => N431);
   C3048 : GTECH_AND2 port map( A => N304, B => plane2_2_25_port, Z => N432);
   C3049 : GTECH_AND2 port map( A => N305, B => plane2_2_24_port, Z => N433);
   C3050 : GTECH_AND2 port map( A => N306, B => plane2_2_23_port, Z => N434);
   C3051 : GTECH_AND2 port map( A => N307, B => plane2_2_22_port, Z => N435);
   C3052 : GTECH_AND2 port map( A => N308, B => plane2_2_21_port, Z => N436);
   C3053 : GTECH_XOR2 port map( A => plane0_2_127_port, B => N309, Z => 
                           perm_output(127));
   C3054 : GTECH_XOR2 port map( A => plane0_2_126_port, B => N310, Z => 
                           perm_output(126));
   C3055 : GTECH_XOR2 port map( A => plane0_2_125_port, B => N311, Z => 
                           perm_output(125));
   C3056 : GTECH_XOR2 port map( A => plane0_2_124_port, B => N312, Z => 
                           perm_output(124));
   C3057 : GTECH_XOR2 port map( A => plane0_2_123_port, B => N313, Z => 
                           perm_output(123));
   C3058 : GTECH_XOR2 port map( A => plane0_2_122_port, B => N314, Z => 
                           perm_output(122));
   C3059 : GTECH_XOR2 port map( A => plane0_2_121_port, B => N315, Z => 
                           perm_output(121));
   C3060 : GTECH_XOR2 port map( A => plane0_2_120_port, B => N316, Z => 
                           perm_output(120));
   C3061 : GTECH_XOR2 port map( A => plane0_2_119_port, B => N317, Z => 
                           perm_output(119));
   C3062 : GTECH_XOR2 port map( A => plane0_2_118_port, B => N318, Z => 
                           perm_output(118));
   C3063 : GTECH_XOR2 port map( A => plane0_2_117_port, B => N319, Z => 
                           perm_output(117));
   C3064 : GTECH_XOR2 port map( A => plane0_2_116_port, B => N320, Z => 
                           perm_output(116));
   C3065 : GTECH_XOR2 port map( A => plane0_2_115_port, B => N321, Z => 
                           perm_output(115));
   C3066 : GTECH_XOR2 port map( A => plane0_2_114_port, B => N322, Z => 
                           perm_output(114));
   C3067 : GTECH_XOR2 port map( A => plane0_2_113_port, B => N323, Z => 
                           perm_output(113));
   C3068 : GTECH_XOR2 port map( A => plane0_2_112_port, B => N324, Z => 
                           perm_output(112));
   C3069 : GTECH_XOR2 port map( A => plane0_2_111_port, B => N325, Z => 
                           perm_output(111));
   C3070 : GTECH_XOR2 port map( A => plane0_2_110_port, B => N326, Z => 
                           perm_output(110));
   C3071 : GTECH_XOR2 port map( A => plane0_2_109_port, B => N327, Z => 
                           perm_output(109));
   C3072 : GTECH_XOR2 port map( A => plane0_2_108_port, B => N328, Z => 
                           perm_output(108));
   C3073 : GTECH_XOR2 port map( A => add_rnd_const_small_11_port, B => N329, Z 
                           => perm_output(107));
   C3074 : GTECH_XOR2 port map( A => add_rnd_const_small_10_port, B => N330, Z 
                           => perm_output(106));
   C3075 : GTECH_XOR2 port map( A => add_rnd_const_small_9_port, B => N331, Z 
                           => perm_output(105));
   C3076 : GTECH_XOR2 port map( A => add_rnd_const_small_8_port, B => N332, Z 
                           => perm_output(104));
   C3077 : GTECH_XOR2 port map( A => add_rnd_const_small_7_port, B => N333, Z 
                           => perm_output(103));
   C3078 : GTECH_XOR2 port map( A => add_rnd_const_small_6_port, B => N334, Z 
                           => perm_output(102));
   C3079 : GTECH_XOR2 port map( A => add_rnd_const_small_5_port, B => N335, Z 
                           => perm_output(101));
   C3080 : GTECH_XOR2 port map( A => add_rnd_const_small_4_port, B => N336, Z 
                           => perm_output(100));
   C3081 : GTECH_XOR2 port map( A => add_rnd_const_small_3_port, B => N337, Z 
                           => perm_output(99));
   C3082 : GTECH_XOR2 port map( A => add_rnd_const_small_2_port, B => N338, Z 
                           => perm_output(98));
   C3083 : GTECH_XOR2 port map( A => add_rnd_const_small_1_port, B => N339, Z 
                           => perm_output(97));
   C3084 : GTECH_XOR2 port map( A => add_rnd_const_small_0_port, B => N340, Z 
                           => perm_output(96));
   C3085 : GTECH_XOR2 port map( A => plane0_2_95_port, B => N341, Z => 
                           perm_output(95));
   C3086 : GTECH_XOR2 port map( A => plane0_2_94_port, B => N342, Z => 
                           perm_output(94));
   C3087 : GTECH_XOR2 port map( A => plane0_2_93_port, B => N343, Z => 
                           perm_output(93));
   C3088 : GTECH_XOR2 port map( A => plane0_2_92_port, B => N344, Z => 
                           perm_output(92));
   C3089 : GTECH_XOR2 port map( A => plane0_2_91_port, B => N345, Z => 
                           perm_output(91));
   C3090 : GTECH_XOR2 port map( A => plane0_2_90_port, B => N346, Z => 
                           perm_output(90));
   C3091 : GTECH_XOR2 port map( A => plane0_2_89_port, B => N347, Z => 
                           perm_output(89));
   C3092 : GTECH_XOR2 port map( A => plane0_2_88_port, B => N348, Z => 
                           perm_output(88));
   C3093 : GTECH_XOR2 port map( A => plane0_2_87_port, B => N349, Z => 
                           perm_output(87));
   C3094 : GTECH_XOR2 port map( A => plane0_2_86_port, B => N350, Z => 
                           perm_output(86));
   C3095 : GTECH_XOR2 port map( A => plane0_2_85_port, B => N351, Z => 
                           perm_output(85));
   C3096 : GTECH_XOR2 port map( A => plane0_2_84_port, B => N352, Z => 
                           perm_output(84));
   C3097 : GTECH_XOR2 port map( A => plane0_2_83_port, B => N353, Z => 
                           perm_output(83));
   C3098 : GTECH_XOR2 port map( A => plane0_2_82_port, B => N354, Z => 
                           perm_output(82));
   C3099 : GTECH_XOR2 port map( A => plane0_2_81_port, B => N355, Z => 
                           perm_output(81));
   C3100 : GTECH_XOR2 port map( A => plane0_2_80_port, B => N356, Z => 
                           perm_output(80));
   C3101 : GTECH_XOR2 port map( A => plane0_2_79_port, B => N357, Z => 
                           perm_output(79));
   C3102 : GTECH_XOR2 port map( A => plane0_2_78_port, B => N358, Z => 
                           perm_output(78));
   C3103 : GTECH_XOR2 port map( A => plane0_2_77_port, B => N359, Z => 
                           perm_output(77));
   C3104 : GTECH_XOR2 port map( A => plane0_2_76_port, B => N360, Z => 
                           perm_output(76));
   C3105 : GTECH_XOR2 port map( A => plane0_2_75_port, B => N361, Z => 
                           perm_output(75));
   C3106 : GTECH_XOR2 port map( A => plane0_2_74_port, B => N362, Z => 
                           perm_output(74));
   C3107 : GTECH_XOR2 port map( A => plane0_2_73_port, B => N363, Z => 
                           perm_output(73));
   C3108 : GTECH_XOR2 port map( A => plane0_2_72_port, B => N364, Z => 
                           perm_output(72));
   C3109 : GTECH_XOR2 port map( A => plane0_2_71_port, B => N365, Z => 
                           perm_output(71));
   C3110 : GTECH_XOR2 port map( A => plane0_2_70_port, B => N366, Z => 
                           perm_output(70));
   C3111 : GTECH_XOR2 port map( A => plane0_2_69_port, B => N367, Z => 
                           perm_output(69));
   C3112 : GTECH_XOR2 port map( A => plane0_2_68_port, B => N368, Z => 
                           perm_output(68));
   C3113 : GTECH_XOR2 port map( A => plane0_2_67_port, B => N369, Z => 
                           perm_output(67));
   C3114 : GTECH_XOR2 port map( A => plane0_2_66_port, B => N370, Z => 
                           perm_output(66));
   C3115 : GTECH_XOR2 port map( A => plane0_2_65_port, B => N371, Z => 
                           perm_output(65));
   C3116 : GTECH_XOR2 port map( A => plane0_2_64_port, B => N372, Z => 
                           perm_output(64));
   C3117 : GTECH_XOR2 port map( A => plane0_2_63_port, B => N373, Z => 
                           perm_output(63));
   C3118 : GTECH_XOR2 port map( A => plane0_2_62_port, B => N374, Z => 
                           perm_output(62));
   C3119 : GTECH_XOR2 port map( A => plane0_2_61_port, B => N375, Z => 
                           perm_output(61));
   C3120 : GTECH_XOR2 port map( A => plane0_2_60_port, B => N376, Z => 
                           perm_output(60));
   C3121 : GTECH_XOR2 port map( A => plane0_2_59_port, B => N377, Z => 
                           perm_output(59));
   C3122 : GTECH_XOR2 port map( A => plane0_2_58_port, B => N378, Z => 
                           perm_output(58));
   C3123 : GTECH_XOR2 port map( A => plane0_2_57_port, B => N379, Z => 
                           perm_output(57));
   C3124 : GTECH_XOR2 port map( A => plane0_2_56_port, B => N380, Z => 
                           perm_output(56));
   C3125 : GTECH_XOR2 port map( A => plane0_2_55_port, B => N381, Z => 
                           perm_output(55));
   C3126 : GTECH_XOR2 port map( A => plane0_2_54_port, B => N382, Z => 
                           perm_output(54));
   C3127 : GTECH_XOR2 port map( A => plane0_2_53_port, B => N383, Z => 
                           perm_output(53));
   C3128 : GTECH_XOR2 port map( A => plane0_2_52_port, B => N384, Z => 
                           perm_output(52));
   C3129 : GTECH_XOR2 port map( A => plane0_2_51_port, B => N385, Z => 
                           perm_output(51));
   C3130 : GTECH_XOR2 port map( A => plane0_2_50_port, B => N386, Z => 
                           perm_output(50));
   C3131 : GTECH_XOR2 port map( A => plane0_2_49_port, B => N387, Z => 
                           perm_output(49));
   C3132 : GTECH_XOR2 port map( A => plane0_2_48_port, B => N388, Z => 
                           perm_output(48));
   C3133 : GTECH_XOR2 port map( A => plane0_2_47_port, B => N389, Z => 
                           perm_output(47));
   C3134 : GTECH_XOR2 port map( A => plane0_2_46_port, B => N390, Z => 
                           perm_output(46));
   C3135 : GTECH_XOR2 port map( A => plane0_2_45_port, B => N391, Z => 
                           perm_output(45));
   C3136 : GTECH_XOR2 port map( A => plane0_2_44_port, B => N392, Z => 
                           perm_output(44));
   C3137 : GTECH_XOR2 port map( A => plane0_2_43_port, B => N393, Z => 
                           perm_output(43));
   C3138 : GTECH_XOR2 port map( A => plane0_2_42_port, B => N394, Z => 
                           perm_output(42));
   C3139 : GTECH_XOR2 port map( A => plane0_2_41_port, B => N395, Z => 
                           perm_output(41));
   C3140 : GTECH_XOR2 port map( A => plane0_2_40_port, B => N396, Z => 
                           perm_output(40));
   C3141 : GTECH_XOR2 port map( A => plane0_2_39_port, B => N397, Z => 
                           perm_output(39));
   C3142 : GTECH_XOR2 port map( A => plane0_2_38_port, B => N398, Z => 
                           perm_output(38));
   C3143 : GTECH_XOR2 port map( A => plane0_2_37_port, B => N399, Z => 
                           perm_output(37));
   C3144 : GTECH_XOR2 port map( A => plane0_2_36_port, B => N400, Z => 
                           perm_output(36));
   C3145 : GTECH_XOR2 port map( A => plane0_2_35_port, B => N401, Z => 
                           perm_output(35));
   C3146 : GTECH_XOR2 port map( A => plane0_2_34_port, B => N402, Z => 
                           perm_output(34));
   C3147 : GTECH_XOR2 port map( A => plane0_2_33_port, B => N403, Z => 
                           perm_output(33));
   C3148 : GTECH_XOR2 port map( A => plane0_2_32_port, B => N404, Z => 
                           perm_output(32));
   C3149 : GTECH_XOR2 port map( A => plane0_2_31_port, B => N405, Z => 
                           perm_output(31));
   C3150 : GTECH_XOR2 port map( A => plane0_2_30_port, B => N406, Z => 
                           perm_output(30));
   C3151 : GTECH_XOR2 port map( A => plane0_2_29_port, B => N407, Z => 
                           perm_output(29));
   C3152 : GTECH_XOR2 port map( A => plane0_2_28_port, B => N408, Z => 
                           perm_output(28));
   C3153 : GTECH_XOR2 port map( A => plane0_2_27_port, B => N409, Z => 
                           perm_output(27));
   C3154 : GTECH_XOR2 port map( A => plane0_2_26_port, B => N410, Z => 
                           perm_output(26));
   C3155 : GTECH_XOR2 port map( A => plane0_2_25_port, B => N411, Z => 
                           perm_output(25));
   C3156 : GTECH_XOR2 port map( A => plane0_2_24_port, B => N412, Z => 
                           perm_output(24));
   C3157 : GTECH_XOR2 port map( A => plane0_2_23_port, B => N413, Z => 
                           perm_output(23));
   C3158 : GTECH_XOR2 port map( A => plane0_2_22_port, B => N414, Z => 
                           perm_output(22));
   C3159 : GTECH_XOR2 port map( A => plane0_2_21_port, B => N415, Z => 
                           perm_output(21));
   C3160 : GTECH_XOR2 port map( A => plane0_2_20_port, B => N416, Z => 
                           perm_output(20));
   C3161 : GTECH_XOR2 port map( A => plane0_2_19_port, B => N417, Z => 
                           perm_output(19));
   C3162 : GTECH_XOR2 port map( A => plane0_2_18_port, B => N418, Z => 
                           perm_output(18));
   C3163 : GTECH_XOR2 port map( A => plane0_2_17_port, B => N419, Z => 
                           perm_output(17));
   C3164 : GTECH_XOR2 port map( A => plane0_2_16_port, B => N420, Z => 
                           perm_output(16));
   C3165 : GTECH_XOR2 port map( A => plane0_2_15_port, B => N421, Z => 
                           perm_output(15));
   C3166 : GTECH_XOR2 port map( A => plane0_2_14_port, B => N422, Z => 
                           perm_output(14));
   C3167 : GTECH_XOR2 port map( A => plane0_2_13_port, B => N423, Z => 
                           perm_output(13));
   C3168 : GTECH_XOR2 port map( A => plane0_2_12_port, B => N424, Z => 
                           perm_output(12));
   C3169 : GTECH_XOR2 port map( A => plane0_2_11_port, B => N425, Z => 
                           perm_output(11));
   C3170 : GTECH_XOR2 port map( A => plane0_2_10_port, B => N426, Z => 
                           perm_output(10));
   C3171 : GTECH_XOR2 port map( A => plane0_2_9_port, B => N427, Z => 
                           perm_output(9));
   C3172 : GTECH_XOR2 port map( A => plane0_2_8_port, B => N428, Z => 
                           perm_output(8));
   C3173 : GTECH_XOR2 port map( A => plane0_2_7_port, B => N429, Z => 
                           perm_output(7));
   C3174 : GTECH_XOR2 port map( A => plane0_2_6_port, B => N430, Z => 
                           perm_output(6));
   C3175 : GTECH_XOR2 port map( A => plane0_2_5_port, B => N431, Z => 
                           perm_output(5));
   C3176 : GTECH_XOR2 port map( A => plane0_2_4_port, B => N432, Z => 
                           perm_output(4));
   C3177 : GTECH_XOR2 port map( A => plane0_2_3_port, B => N433, Z => 
                           perm_output(3));
   C3178 : GTECH_XOR2 port map( A => plane0_2_2_port, B => N434, Z => 
                           perm_output(2));
   C3179 : GTECH_XOR2 port map( A => plane0_2_1_port, B => N435, Z => 
                           perm_output(1));
   C3180 : GTECH_XOR2 port map( A => plane0_2_0_port, B => N436, Z => 
                           perm_output(0));
   I_148 : GTECH_NOT port map( A => plane2_2_116_port, Z => N437);
   I_149 : GTECH_NOT port map( A => plane2_2_115_port, Z => N438);
   I_150 : GTECH_NOT port map( A => plane2_2_114_port, Z => N439);
   I_151 : GTECH_NOT port map( A => plane2_2_113_port, Z => N440);
   I_152 : GTECH_NOT port map( A => plane2_2_112_port, Z => N441);
   I_153 : GTECH_NOT port map( A => plane2_2_111_port, Z => N442);
   I_154 : GTECH_NOT port map( A => plane2_2_110_port, Z => N443);
   I_155 : GTECH_NOT port map( A => plane2_2_109_port, Z => N444);
   I_156 : GTECH_NOT port map( A => plane2_2_108_port, Z => N445);
   I_157 : GTECH_NOT port map( A => plane2_2_107_port, Z => N446);
   I_158 : GTECH_NOT port map( A => plane2_2_106_port, Z => N447);
   I_159 : GTECH_NOT port map( A => plane2_2_105_port, Z => N448);
   I_160 : GTECH_NOT port map( A => plane2_2_104_port, Z => N449);
   I_161 : GTECH_NOT port map( A => plane2_2_103_port, Z => N450);
   I_162 : GTECH_NOT port map( A => plane2_2_102_port, Z => N451);
   I_163 : GTECH_NOT port map( A => plane2_2_101_port, Z => N452);
   I_164 : GTECH_NOT port map( A => plane2_2_100_port, Z => N453);
   I_165 : GTECH_NOT port map( A => plane2_2_99_port, Z => N454);
   I_166 : GTECH_NOT port map( A => plane2_2_98_port, Z => N455);
   I_167 : GTECH_NOT port map( A => plane2_2_97_port, Z => N456);
   I_168 : GTECH_NOT port map( A => plane2_2_96_port, Z => N457);
   I_169 : GTECH_NOT port map( A => plane2_2_127_port, Z => N458);
   I_170 : GTECH_NOT port map( A => plane2_2_126_port, Z => N459);
   I_171 : GTECH_NOT port map( A => plane2_2_125_port, Z => N460);
   I_172 : GTECH_NOT port map( A => plane2_2_124_port, Z => N461);
   I_173 : GTECH_NOT port map( A => plane2_2_123_port, Z => N462);
   I_174 : GTECH_NOT port map( A => plane2_2_122_port, Z => N463);
   I_175 : GTECH_NOT port map( A => plane2_2_121_port, Z => N464);
   I_176 : GTECH_NOT port map( A => plane2_2_120_port, Z => N465);
   I_177 : GTECH_NOT port map( A => plane2_2_119_port, Z => N466);
   I_178 : GTECH_NOT port map( A => plane2_2_118_port, Z => N467);
   I_179 : GTECH_NOT port map( A => plane2_2_117_port, Z => N468);
   I_180 : GTECH_NOT port map( A => plane2_2_84_port, Z => N469);
   I_181 : GTECH_NOT port map( A => plane2_2_83_port, Z => N470);
   I_182 : GTECH_NOT port map( A => plane2_2_82_port, Z => N471);
   I_183 : GTECH_NOT port map( A => plane2_2_81_port, Z => N472);
   I_184 : GTECH_NOT port map( A => plane2_2_80_port, Z => N473);
   I_185 : GTECH_NOT port map( A => plane2_2_79_port, Z => N474);
   I_186 : GTECH_NOT port map( A => plane2_2_78_port, Z => N475);
   I_187 : GTECH_NOT port map( A => plane2_2_77_port, Z => N476);
   I_188 : GTECH_NOT port map( A => plane2_2_76_port, Z => N477);
   I_189 : GTECH_NOT port map( A => plane2_2_75_port, Z => N478);
   I_190 : GTECH_NOT port map( A => plane2_2_74_port, Z => N479);
   I_191 : GTECH_NOT port map( A => plane2_2_73_port, Z => N480);
   I_192 : GTECH_NOT port map( A => plane2_2_72_port, Z => N481);
   I_193 : GTECH_NOT port map( A => plane2_2_71_port, Z => N482);
   I_194 : GTECH_NOT port map( A => plane2_2_70_port, Z => N483);
   I_195 : GTECH_NOT port map( A => plane2_2_69_port, Z => N484);
   I_196 : GTECH_NOT port map( A => plane2_2_68_port, Z => N485);
   I_197 : GTECH_NOT port map( A => plane2_2_67_port, Z => N486);
   I_198 : GTECH_NOT port map( A => plane2_2_66_port, Z => N487);
   I_199 : GTECH_NOT port map( A => plane2_2_65_port, Z => N488);
   I_200 : GTECH_NOT port map( A => plane2_2_64_port, Z => N489);
   I_201 : GTECH_NOT port map( A => plane2_2_95_port, Z => N490);
   I_202 : GTECH_NOT port map( A => plane2_2_94_port, Z => N491);
   I_203 : GTECH_NOT port map( A => plane2_2_93_port, Z => N492);
   I_204 : GTECH_NOT port map( A => plane2_2_92_port, Z => N493);
   I_205 : GTECH_NOT port map( A => plane2_2_91_port, Z => N494);
   I_206 : GTECH_NOT port map( A => plane2_2_90_port, Z => N495);
   I_207 : GTECH_NOT port map( A => plane2_2_89_port, Z => N496);
   I_208 : GTECH_NOT port map( A => plane2_2_88_port, Z => N497);
   I_209 : GTECH_NOT port map( A => plane2_2_87_port, Z => N498);
   I_210 : GTECH_NOT port map( A => plane2_2_86_port, Z => N499);
   I_211 : GTECH_NOT port map( A => plane2_2_85_port, Z => N500);
   I_212 : GTECH_NOT port map( A => plane2_2_52_port, Z => N501);
   I_213 : GTECH_NOT port map( A => plane2_2_51_port, Z => N502);
   I_214 : GTECH_NOT port map( A => plane2_2_50_port, Z => N503);
   I_215 : GTECH_NOT port map( A => plane2_2_49_port, Z => N504);
   I_216 : GTECH_NOT port map( A => plane2_2_48_port, Z => N505);
   I_217 : GTECH_NOT port map( A => plane2_2_47_port, Z => N506);
   I_218 : GTECH_NOT port map( A => plane2_2_46_port, Z => N507);
   I_219 : GTECH_NOT port map( A => plane2_2_45_port, Z => N508);
   I_220 : GTECH_NOT port map( A => plane2_2_44_port, Z => N509);
   I_221 : GTECH_NOT port map( A => plane2_2_43_port, Z => N510);
   I_222 : GTECH_NOT port map( A => plane2_2_42_port, Z => N511);
   I_223 : GTECH_NOT port map( A => plane2_2_41_port, Z => N512);
   I_224 : GTECH_NOT port map( A => plane2_2_40_port, Z => N513);
   I_225 : GTECH_NOT port map( A => plane2_2_39_port, Z => N514);
   I_226 : GTECH_NOT port map( A => plane2_2_38_port, Z => N515);
   I_227 : GTECH_NOT port map( A => plane2_2_37_port, Z => N516);
   I_228 : GTECH_NOT port map( A => plane2_2_36_port, Z => N517);
   I_229 : GTECH_NOT port map( A => plane2_2_35_port, Z => N518);
   I_230 : GTECH_NOT port map( A => plane2_2_34_port, Z => N519);
   I_231 : GTECH_NOT port map( A => plane2_2_33_port, Z => N520);
   I_232 : GTECH_NOT port map( A => plane2_2_32_port, Z => N521);
   I_233 : GTECH_NOT port map( A => plane2_2_63_port, Z => N522);
   I_234 : GTECH_NOT port map( A => plane2_2_62_port, Z => N523);
   I_235 : GTECH_NOT port map( A => plane2_2_61_port, Z => N524);
   I_236 : GTECH_NOT port map( A => plane2_2_60_port, Z => N525);
   I_237 : GTECH_NOT port map( A => plane2_2_59_port, Z => N526);
   I_238 : GTECH_NOT port map( A => plane2_2_58_port, Z => N527);
   I_239 : GTECH_NOT port map( A => plane2_2_57_port, Z => N528);
   I_240 : GTECH_NOT port map( A => plane2_2_56_port, Z => N529);
   I_241 : GTECH_NOT port map( A => plane2_2_55_port, Z => N530);
   I_242 : GTECH_NOT port map( A => plane2_2_54_port, Z => N531);
   I_243 : GTECH_NOT port map( A => plane2_2_53_port, Z => N532);
   I_244 : GTECH_NOT port map( A => plane2_2_20_port, Z => N533);
   I_245 : GTECH_NOT port map( A => plane2_2_19_port, Z => N534);
   I_246 : GTECH_NOT port map( A => plane2_2_18_port, Z => N535);
   I_247 : GTECH_NOT port map( A => plane2_2_17_port, Z => N536);
   I_248 : GTECH_NOT port map( A => plane2_2_16_port, Z => N537);
   I_249 : GTECH_NOT port map( A => plane2_2_15_port, Z => N538);
   I_250 : GTECH_NOT port map( A => plane2_2_14_port, Z => N539);
   I_251 : GTECH_NOT port map( A => plane2_2_13_port, Z => N540);
   I_252 : GTECH_NOT port map( A => plane2_2_12_port, Z => N541);
   I_253 : GTECH_NOT port map( A => plane2_2_11_port, Z => N542);
   I_254 : GTECH_NOT port map( A => plane2_2_10_port, Z => N543);
   I_255 : GTECH_NOT port map( A => plane2_2_9_port, Z => N544);
   I_256 : GTECH_NOT port map( A => plane2_2_8_port, Z => N545);
   I_257 : GTECH_NOT port map( A => plane2_2_7_port, Z => N546);
   I_258 : GTECH_NOT port map( A => plane2_2_6_port, Z => N547);
   I_259 : GTECH_NOT port map( A => plane2_2_5_port, Z => N548);
   I_260 : GTECH_NOT port map( A => plane2_2_4_port, Z => N549);
   I_261 : GTECH_NOT port map( A => plane2_2_3_port, Z => N550);
   I_262 : GTECH_NOT port map( A => plane2_2_2_port, Z => N551);
   I_263 : GTECH_NOT port map( A => plane2_2_1_port, Z => N552);
   I_264 : GTECH_NOT port map( A => plane2_2_0_port, Z => N553);
   I_265 : GTECH_NOT port map( A => plane2_2_31_port, Z => N554);
   I_266 : GTECH_NOT port map( A => plane2_2_30_port, Z => N555);
   I_267 : GTECH_NOT port map( A => plane2_2_29_port, Z => N556);
   I_268 : GTECH_NOT port map( A => plane2_2_28_port, Z => N557);
   I_269 : GTECH_NOT port map( A => plane2_2_27_port, Z => N558);
   I_270 : GTECH_NOT port map( A => plane2_2_26_port, Z => N559);
   I_271 : GTECH_NOT port map( A => plane2_2_25_port, Z => N560);
   I_272 : GTECH_NOT port map( A => plane2_2_24_port, Z => N561);
   I_273 : GTECH_NOT port map( A => plane2_2_23_port, Z => N562);
   I_274 : GTECH_NOT port map( A => plane2_2_22_port, Z => N563);
   I_275 : GTECH_NOT port map( A => plane2_2_21_port, Z => N564);
   C3309 : GTECH_AND2 port map( A => N437, B => plane0_2_127_port, Z => N565);
   C3310 : GTECH_AND2 port map( A => N438, B => plane0_2_126_port, Z => N566);
   C3311 : GTECH_AND2 port map( A => N439, B => plane0_2_125_port, Z => N567);
   C3312 : GTECH_AND2 port map( A => N440, B => plane0_2_124_port, Z => N568);
   C3313 : GTECH_AND2 port map( A => N441, B => plane0_2_123_port, Z => N569);
   C3314 : GTECH_AND2 port map( A => N442, B => plane0_2_122_port, Z => N570);
   C3315 : GTECH_AND2 port map( A => N443, B => plane0_2_121_port, Z => N571);
   C3316 : GTECH_AND2 port map( A => N444, B => plane0_2_120_port, Z => N572);
   C3317 : GTECH_AND2 port map( A => N445, B => plane0_2_119_port, Z => N573);
   C3318 : GTECH_AND2 port map( A => N446, B => plane0_2_118_port, Z => N574);
   C3319 : GTECH_AND2 port map( A => N447, B => plane0_2_117_port, Z => N575);
   C3320 : GTECH_AND2 port map( A => N448, B => plane0_2_116_port, Z => N576);
   C3321 : GTECH_AND2 port map( A => N449, B => plane0_2_115_port, Z => N577);
   C3322 : GTECH_AND2 port map( A => N450, B => plane0_2_114_port, Z => N578);
   C3323 : GTECH_AND2 port map( A => N451, B => plane0_2_113_port, Z => N579);
   C3324 : GTECH_AND2 port map( A => N452, B => plane0_2_112_port, Z => N580);
   C3325 : GTECH_AND2 port map( A => N453, B => plane0_2_111_port, Z => N581);
   C3326 : GTECH_AND2 port map( A => N454, B => plane0_2_110_port, Z => N582);
   C3327 : GTECH_AND2 port map( A => N455, B => plane0_2_109_port, Z => N583);
   C3328 : GTECH_AND2 port map( A => N456, B => plane0_2_108_port, Z => N584);
   C3329 : GTECH_AND2 port map( A => N457, B => add_rnd_const_small_11_port, Z 
                           => N585);
   C3330 : GTECH_AND2 port map( A => N458, B => add_rnd_const_small_10_port, Z 
                           => N586);
   C3331 : GTECH_AND2 port map( A => N459, B => add_rnd_const_small_9_port, Z 
                           => N587);
   C3332 : GTECH_AND2 port map( A => N460, B => add_rnd_const_small_8_port, Z 
                           => N588);
   C3333 : GTECH_AND2 port map( A => N461, B => add_rnd_const_small_7_port, Z 
                           => N589);
   C3334 : GTECH_AND2 port map( A => N462, B => add_rnd_const_small_6_port, Z 
                           => N590);
   C3335 : GTECH_AND2 port map( A => N463, B => add_rnd_const_small_5_port, Z 
                           => N591);
   C3336 : GTECH_AND2 port map( A => N464, B => add_rnd_const_small_4_port, Z 
                           => N592);
   C3337 : GTECH_AND2 port map( A => N465, B => add_rnd_const_small_3_port, Z 
                           => N593);
   C3338 : GTECH_AND2 port map( A => N466, B => add_rnd_const_small_2_port, Z 
                           => N594);
   C3339 : GTECH_AND2 port map( A => N467, B => add_rnd_const_small_1_port, Z 
                           => N595);
   C3340 : GTECH_AND2 port map( A => N468, B => add_rnd_const_small_0_port, Z 
                           => N596);
   C3341 : GTECH_AND2 port map( A => N469, B => plane0_2_95_port, Z => N597);
   C3342 : GTECH_AND2 port map( A => N470, B => plane0_2_94_port, Z => N598);
   C3343 : GTECH_AND2 port map( A => N471, B => plane0_2_93_port, Z => N599);
   C3344 : GTECH_AND2 port map( A => N472, B => plane0_2_92_port, Z => N600);
   C3345 : GTECH_AND2 port map( A => N473, B => plane0_2_91_port, Z => N601);
   C3346 : GTECH_AND2 port map( A => N474, B => plane0_2_90_port, Z => N602);
   C3347 : GTECH_AND2 port map( A => N475, B => plane0_2_89_port, Z => N603);
   C3348 : GTECH_AND2 port map( A => N476, B => plane0_2_88_port, Z => N604);
   C3349 : GTECH_AND2 port map( A => N477, B => plane0_2_87_port, Z => N605);
   C3350 : GTECH_AND2 port map( A => N478, B => plane0_2_86_port, Z => N606);
   C3351 : GTECH_AND2 port map( A => N479, B => plane0_2_85_port, Z => N607);
   C3352 : GTECH_AND2 port map( A => N480, B => plane0_2_84_port, Z => N608);
   C3353 : GTECH_AND2 port map( A => N481, B => plane0_2_83_port, Z => N609);
   C3354 : GTECH_AND2 port map( A => N482, B => plane0_2_82_port, Z => N610);
   C3355 : GTECH_AND2 port map( A => N483, B => plane0_2_81_port, Z => N611);
   C3356 : GTECH_AND2 port map( A => N484, B => plane0_2_80_port, Z => N612);
   C3357 : GTECH_AND2 port map( A => N485, B => plane0_2_79_port, Z => N613);
   C3358 : GTECH_AND2 port map( A => N486, B => plane0_2_78_port, Z => N614);
   C3359 : GTECH_AND2 port map( A => N487, B => plane0_2_77_port, Z => N615);
   C3360 : GTECH_AND2 port map( A => N488, B => plane0_2_76_port, Z => N616);
   C3361 : GTECH_AND2 port map( A => N489, B => plane0_2_75_port, Z => N617);
   C3362 : GTECH_AND2 port map( A => N490, B => plane0_2_74_port, Z => N618);
   C3363 : GTECH_AND2 port map( A => N491, B => plane0_2_73_port, Z => N619);
   C3364 : GTECH_AND2 port map( A => N492, B => plane0_2_72_port, Z => N620);
   C3365 : GTECH_AND2 port map( A => N493, B => plane0_2_71_port, Z => N621);
   C3366 : GTECH_AND2 port map( A => N494, B => plane0_2_70_port, Z => N622);
   C3367 : GTECH_AND2 port map( A => N495, B => plane0_2_69_port, Z => N623);
   C3368 : GTECH_AND2 port map( A => N496, B => plane0_2_68_port, Z => N624);
   C3369 : GTECH_AND2 port map( A => N497, B => plane0_2_67_port, Z => N625);
   C3370 : GTECH_AND2 port map( A => N498, B => plane0_2_66_port, Z => N626);
   C3371 : GTECH_AND2 port map( A => N499, B => plane0_2_65_port, Z => N627);
   C3372 : GTECH_AND2 port map( A => N500, B => plane0_2_64_port, Z => N628);
   C3373 : GTECH_AND2 port map( A => N501, B => plane0_2_63_port, Z => N629);
   C3374 : GTECH_AND2 port map( A => N502, B => plane0_2_62_port, Z => N630);
   C3375 : GTECH_AND2 port map( A => N503, B => plane0_2_61_port, Z => N631);
   C3376 : GTECH_AND2 port map( A => N504, B => plane0_2_60_port, Z => N632);
   C3377 : GTECH_AND2 port map( A => N505, B => plane0_2_59_port, Z => N633);
   C3378 : GTECH_AND2 port map( A => N506, B => plane0_2_58_port, Z => N634);
   C3379 : GTECH_AND2 port map( A => N507, B => plane0_2_57_port, Z => N635);
   C3380 : GTECH_AND2 port map( A => N508, B => plane0_2_56_port, Z => N636);
   C3381 : GTECH_AND2 port map( A => N509, B => plane0_2_55_port, Z => N637);
   C3382 : GTECH_AND2 port map( A => N510, B => plane0_2_54_port, Z => N638);
   C3383 : GTECH_AND2 port map( A => N511, B => plane0_2_53_port, Z => N639);
   C3384 : GTECH_AND2 port map( A => N512, B => plane0_2_52_port, Z => N640);
   C3385 : GTECH_AND2 port map( A => N513, B => plane0_2_51_port, Z => N641);
   C3386 : GTECH_AND2 port map( A => N514, B => plane0_2_50_port, Z => N642);
   C3387 : GTECH_AND2 port map( A => N515, B => plane0_2_49_port, Z => N643);
   C3388 : GTECH_AND2 port map( A => N516, B => plane0_2_48_port, Z => N644);
   C3389 : GTECH_AND2 port map( A => N517, B => plane0_2_47_port, Z => N645);
   C3390 : GTECH_AND2 port map( A => N518, B => plane0_2_46_port, Z => N646);
   C3391 : GTECH_AND2 port map( A => N519, B => plane0_2_45_port, Z => N647);
   C3392 : GTECH_AND2 port map( A => N520, B => plane0_2_44_port, Z => N648);
   C3393 : GTECH_AND2 port map( A => N521, B => plane0_2_43_port, Z => N649);
   C3394 : GTECH_AND2 port map( A => N522, B => plane0_2_42_port, Z => N650);
   C3395 : GTECH_AND2 port map( A => N523, B => plane0_2_41_port, Z => N651);
   C3396 : GTECH_AND2 port map( A => N524, B => plane0_2_40_port, Z => N652);
   C3397 : GTECH_AND2 port map( A => N525, B => plane0_2_39_port, Z => N653);
   C3398 : GTECH_AND2 port map( A => N526, B => plane0_2_38_port, Z => N654);
   C3399 : GTECH_AND2 port map( A => N527, B => plane0_2_37_port, Z => N655);
   C3400 : GTECH_AND2 port map( A => N528, B => plane0_2_36_port, Z => N656);
   C3401 : GTECH_AND2 port map( A => N529, B => plane0_2_35_port, Z => N657);
   C3402 : GTECH_AND2 port map( A => N530, B => plane0_2_34_port, Z => N658);
   C3403 : GTECH_AND2 port map( A => N531, B => plane0_2_33_port, Z => N659);
   C3404 : GTECH_AND2 port map( A => N532, B => plane0_2_32_port, Z => N660);
   C3405 : GTECH_AND2 port map( A => N533, B => plane0_2_31_port, Z => N661);
   C3406 : GTECH_AND2 port map( A => N534, B => plane0_2_30_port, Z => N662);
   C3407 : GTECH_AND2 port map( A => N535, B => plane0_2_29_port, Z => N663);
   C3408 : GTECH_AND2 port map( A => N536, B => plane0_2_28_port, Z => N664);
   C3409 : GTECH_AND2 port map( A => N537, B => plane0_2_27_port, Z => N665);
   C3410 : GTECH_AND2 port map( A => N538, B => plane0_2_26_port, Z => N666);
   C3411 : GTECH_AND2 port map( A => N539, B => plane0_2_25_port, Z => N667);
   C3412 : GTECH_AND2 port map( A => N540, B => plane0_2_24_port, Z => N668);
   C3413 : GTECH_AND2 port map( A => N541, B => plane0_2_23_port, Z => N669);
   C3414 : GTECH_AND2 port map( A => N542, B => plane0_2_22_port, Z => N670);
   C3415 : GTECH_AND2 port map( A => N543, B => plane0_2_21_port, Z => N671);
   C3416 : GTECH_AND2 port map( A => N544, B => plane0_2_20_port, Z => N672);
   C3417 : GTECH_AND2 port map( A => N545, B => plane0_2_19_port, Z => N673);
   C3418 : GTECH_AND2 port map( A => N546, B => plane0_2_18_port, Z => N674);
   C3419 : GTECH_AND2 port map( A => N547, B => plane0_2_17_port, Z => N675);
   C3420 : GTECH_AND2 port map( A => N548, B => plane0_2_16_port, Z => N676);
   C3421 : GTECH_AND2 port map( A => N549, B => plane0_2_15_port, Z => N677);
   C3422 : GTECH_AND2 port map( A => N550, B => plane0_2_14_port, Z => N678);
   C3423 : GTECH_AND2 port map( A => N551, B => plane0_2_13_port, Z => N679);
   C3424 : GTECH_AND2 port map( A => N552, B => plane0_2_12_port, Z => N680);
   C3425 : GTECH_AND2 port map( A => N553, B => plane0_2_11_port, Z => N681);
   C3426 : GTECH_AND2 port map( A => N554, B => plane0_2_10_port, Z => N682);
   C3427 : GTECH_AND2 port map( A => N555, B => plane0_2_9_port, Z => N683);
   C3428 : GTECH_AND2 port map( A => N556, B => plane0_2_8_port, Z => N684);
   C3429 : GTECH_AND2 port map( A => N557, B => plane0_2_7_port, Z => N685);
   C3430 : GTECH_AND2 port map( A => N558, B => plane0_2_6_port, Z => N686);
   C3431 : GTECH_AND2 port map( A => N559, B => plane0_2_5_port, Z => N687);
   C3432 : GTECH_AND2 port map( A => N560, B => plane0_2_4_port, Z => N688);
   C3433 : GTECH_AND2 port map( A => N561, B => plane0_2_3_port, Z => N689);
   C3434 : GTECH_AND2 port map( A => N562, B => plane0_2_2_port, Z => N690);
   C3435 : GTECH_AND2 port map( A => N563, B => plane0_2_1_port, Z => N691);
   C3436 : GTECH_AND2 port map( A => N564, B => plane0_2_0_port, Z => N692);
   C3437 : GTECH_XOR2 port map( A => plane1_2_31_port, B => N565, Z => 
                           perm_output(224));
   C3438 : GTECH_XOR2 port map( A => plane1_2_30_port, B => N566, Z => 
                           perm_output(255));
   C3439 : GTECH_XOR2 port map( A => plane1_2_29_port, B => N567, Z => 
                           perm_output(254));
   C3440 : GTECH_XOR2 port map( A => plane1_2_28_port, B => N568, Z => 
                           perm_output(253));
   C3441 : GTECH_XOR2 port map( A => plane1_2_27_port, B => N569, Z => 
                           perm_output(252));
   C3442 : GTECH_XOR2 port map( A => plane1_2_26_port, B => N570, Z => 
                           perm_output(251));
   C3443 : GTECH_XOR2 port map( A => plane1_2_25_port, B => N571, Z => 
                           perm_output(250));
   C3444 : GTECH_XOR2 port map( A => plane1_2_24_port, B => N572, Z => 
                           perm_output(249));
   C3445 : GTECH_XOR2 port map( A => plane1_2_23_port, B => N573, Z => 
                           perm_output(248));
   C3446 : GTECH_XOR2 port map( A => plane1_2_22_port, B => N574, Z => 
                           perm_output(247));
   C3447 : GTECH_XOR2 port map( A => plane1_2_21_port, B => N575, Z => 
                           perm_output(246));
   C3448 : GTECH_XOR2 port map( A => plane1_2_20_port, B => N576, Z => 
                           perm_output(245));
   C3449 : GTECH_XOR2 port map( A => plane1_2_19_port, B => N577, Z => 
                           perm_output(244));
   C3450 : GTECH_XOR2 port map( A => plane1_2_18_port, B => N578, Z => 
                           perm_output(243));
   C3451 : GTECH_XOR2 port map( A => plane1_2_17_port, B => N579, Z => 
                           perm_output(242));
   C3452 : GTECH_XOR2 port map( A => plane1_2_16_port, B => N580, Z => 
                           perm_output(241));
   C3453 : GTECH_XOR2 port map( A => plane1_2_15_port, B => N581, Z => 
                           perm_output(240));
   C3454 : GTECH_XOR2 port map( A => plane1_2_14_port, B => N582, Z => 
                           perm_output(239));
   C3455 : GTECH_XOR2 port map( A => plane1_2_13_port, B => N583, Z => 
                           perm_output(238));
   C3456 : GTECH_XOR2 port map( A => plane1_2_12_port, B => N584, Z => 
                           perm_output(237));
   C3457 : GTECH_XOR2 port map( A => plane1_2_11_port, B => N585, Z => 
                           perm_output(236));
   C3458 : GTECH_XOR2 port map( A => plane1_2_10_port, B => N586, Z => 
                           perm_output(235));
   C3459 : GTECH_XOR2 port map( A => plane1_2_9_port, B => N587, Z => 
                           perm_output(234));
   C3460 : GTECH_XOR2 port map( A => plane1_2_8_port, B => N588, Z => 
                           perm_output(233));
   C3461 : GTECH_XOR2 port map( A => plane1_2_7_port, B => N589, Z => 
                           perm_output(232));
   C3462 : GTECH_XOR2 port map( A => plane1_2_6_port, B => N590, Z => 
                           perm_output(231));
   C3463 : GTECH_XOR2 port map( A => plane1_2_5_port, B => N591, Z => 
                           perm_output(230));
   C3464 : GTECH_XOR2 port map( A => plane1_2_4_port, B => N592, Z => 
                           perm_output(229));
   C3465 : GTECH_XOR2 port map( A => plane1_2_3_port, B => N593, Z => 
                           perm_output(228));
   C3466 : GTECH_XOR2 port map( A => plane1_2_2_port, B => N594, Z => 
                           perm_output(227));
   C3467 : GTECH_XOR2 port map( A => plane1_2_1_port, B => N595, Z => 
                           perm_output(226));
   C3468 : GTECH_XOR2 port map( A => plane1_2_0_port, B => N596, Z => 
                           perm_output(225));
   C3469 : GTECH_XOR2 port map( A => plane1_2_127_port, B => N597, Z => 
                           perm_output(192));
   C3470 : GTECH_XOR2 port map( A => plane1_2_126_port, B => N598, Z => 
                           perm_output(223));
   C3471 : GTECH_XOR2 port map( A => plane1_2_125_port, B => N599, Z => 
                           perm_output(222));
   C3472 : GTECH_XOR2 port map( A => plane1_2_124_port, B => N600, Z => 
                           perm_output(221));
   C3473 : GTECH_XOR2 port map( A => plane1_2_123_port, B => N601, Z => 
                           perm_output(220));
   C3474 : GTECH_XOR2 port map( A => plane1_2_122_port, B => N602, Z => 
                           perm_output(219));
   C3475 : GTECH_XOR2 port map( A => plane1_2_121_port, B => N603, Z => 
                           perm_output(218));
   C3476 : GTECH_XOR2 port map( A => plane1_2_120_port, B => N604, Z => 
                           perm_output(217));
   C3477 : GTECH_XOR2 port map( A => plane1_2_119_port, B => N605, Z => 
                           perm_output(216));
   C3478 : GTECH_XOR2 port map( A => plane1_2_118_port, B => N606, Z => 
                           perm_output(215));
   C3479 : GTECH_XOR2 port map( A => plane1_2_117_port, B => N607, Z => 
                           perm_output(214));
   C3480 : GTECH_XOR2 port map( A => plane1_2_116_port, B => N608, Z => 
                           perm_output(213));
   C3481 : GTECH_XOR2 port map( A => plane1_2_115_port, B => N609, Z => 
                           perm_output(212));
   C3482 : GTECH_XOR2 port map( A => plane1_2_114_port, B => N610, Z => 
                           perm_output(211));
   C3483 : GTECH_XOR2 port map( A => plane1_2_113_port, B => N611, Z => 
                           perm_output(210));
   C3484 : GTECH_XOR2 port map( A => plane1_2_112_port, B => N612, Z => 
                           perm_output(209));
   C3485 : GTECH_XOR2 port map( A => plane1_2_111_port, B => N613, Z => 
                           perm_output(208));
   C3486 : GTECH_XOR2 port map( A => plane1_2_110_port, B => N614, Z => 
                           perm_output(207));
   C3487 : GTECH_XOR2 port map( A => plane1_2_109_port, B => N615, Z => 
                           perm_output(206));
   C3488 : GTECH_XOR2 port map( A => plane1_2_108_port, B => N616, Z => 
                           perm_output(205));
   C3489 : GTECH_XOR2 port map( A => plane1_2_107_port, B => N617, Z => 
                           perm_output(204));
   C3490 : GTECH_XOR2 port map( A => plane1_2_106_port, B => N618, Z => 
                           perm_output(203));
   C3491 : GTECH_XOR2 port map( A => plane1_2_105_port, B => N619, Z => 
                           perm_output(202));
   C3492 : GTECH_XOR2 port map( A => plane1_2_104_port, B => N620, Z => 
                           perm_output(201));
   C3493 : GTECH_XOR2 port map( A => plane1_2_103_port, B => N621, Z => 
                           perm_output(200));
   C3494 : GTECH_XOR2 port map( A => plane1_2_102_port, B => N622, Z => 
                           perm_output(199));
   C3495 : GTECH_XOR2 port map( A => plane1_2_101_port, B => N623, Z => 
                           perm_output(198));
   C3496 : GTECH_XOR2 port map( A => plane1_2_100_port, B => N624, Z => 
                           perm_output(197));
   C3497 : GTECH_XOR2 port map( A => plane1_2_99_port, B => N625, Z => 
                           perm_output(196));
   C3498 : GTECH_XOR2 port map( A => plane1_2_98_port, B => N626, Z => 
                           perm_output(195));
   C3499 : GTECH_XOR2 port map( A => plane1_2_97_port, B => N627, Z => 
                           perm_output(194));
   C3500 : GTECH_XOR2 port map( A => plane1_2_96_port, B => N628, Z => 
                           perm_output(193));
   C3501 : GTECH_XOR2 port map( A => plane1_2_95_port, B => N629, Z => 
                           perm_output(160));
   C3502 : GTECH_XOR2 port map( A => plane1_2_94_port, B => N630, Z => 
                           perm_output(191));
   C3503 : GTECH_XOR2 port map( A => plane1_2_93_port, B => N631, Z => 
                           perm_output(190));
   C3504 : GTECH_XOR2 port map( A => plane1_2_92_port, B => N632, Z => 
                           perm_output(189));
   C3505 : GTECH_XOR2 port map( A => plane1_2_91_port, B => N633, Z => 
                           perm_output(188));
   C3506 : GTECH_XOR2 port map( A => plane1_2_90_port, B => N634, Z => 
                           perm_output(187));
   C3507 : GTECH_XOR2 port map( A => plane1_2_89_port, B => N635, Z => 
                           perm_output(186));
   C3508 : GTECH_XOR2 port map( A => plane1_2_88_port, B => N636, Z => 
                           perm_output(185));
   C3509 : GTECH_XOR2 port map( A => plane1_2_87_port, B => N637, Z => 
                           perm_output(184));
   C3510 : GTECH_XOR2 port map( A => plane1_2_86_port, B => N638, Z => 
                           perm_output(183));
   C3511 : GTECH_XOR2 port map( A => plane1_2_85_port, B => N639, Z => 
                           perm_output(182));
   C3512 : GTECH_XOR2 port map( A => plane1_2_84_port, B => N640, Z => 
                           perm_output(181));
   C3513 : GTECH_XOR2 port map( A => plane1_2_83_port, B => N641, Z => 
                           perm_output(180));
   C3514 : GTECH_XOR2 port map( A => plane1_2_82_port, B => N642, Z => 
                           perm_output(179));
   C3515 : GTECH_XOR2 port map( A => plane1_2_81_port, B => N643, Z => 
                           perm_output(178));
   C3516 : GTECH_XOR2 port map( A => plane1_2_80_port, B => N644, Z => 
                           perm_output(177));
   C3517 : GTECH_XOR2 port map( A => plane1_2_79_port, B => N645, Z => 
                           perm_output(176));
   C3518 : GTECH_XOR2 port map( A => plane1_2_78_port, B => N646, Z => 
                           perm_output(175));
   C3519 : GTECH_XOR2 port map( A => plane1_2_77_port, B => N647, Z => 
                           perm_output(174));
   C3520 : GTECH_XOR2 port map( A => plane1_2_76_port, B => N648, Z => 
                           perm_output(173));
   C3521 : GTECH_XOR2 port map( A => plane1_2_75_port, B => N649, Z => 
                           perm_output(172));
   C3522 : GTECH_XOR2 port map( A => plane1_2_74_port, B => N650, Z => 
                           perm_output(171));
   C3523 : GTECH_XOR2 port map( A => plane1_2_73_port, B => N651, Z => 
                           perm_output(170));
   C3524 : GTECH_XOR2 port map( A => plane1_2_72_port, B => N652, Z => 
                           perm_output(169));
   C3525 : GTECH_XOR2 port map( A => plane1_2_71_port, B => N653, Z => 
                           perm_output(168));
   C3526 : GTECH_XOR2 port map( A => plane1_2_70_port, B => N654, Z => 
                           perm_output(167));
   C3527 : GTECH_XOR2 port map( A => plane1_2_69_port, B => N655, Z => 
                           perm_output(166));
   C3528 : GTECH_XOR2 port map( A => plane1_2_68_port, B => N656, Z => 
                           perm_output(165));
   C3529 : GTECH_XOR2 port map( A => plane1_2_67_port, B => N657, Z => 
                           perm_output(164));
   C3530 : GTECH_XOR2 port map( A => plane1_2_66_port, B => N658, Z => 
                           perm_output(163));
   C3531 : GTECH_XOR2 port map( A => plane1_2_65_port, B => N659, Z => 
                           perm_output(162));
   C3532 : GTECH_XOR2 port map( A => plane1_2_64_port, B => N660, Z => 
                           perm_output(161));
   C3533 : GTECH_XOR2 port map( A => plane1_2_63_port, B => N661, Z => 
                           perm_output(128));
   C3534 : GTECH_XOR2 port map( A => plane1_2_62_port, B => N662, Z => 
                           perm_output(159));
   C3535 : GTECH_XOR2 port map( A => plane1_2_61_port, B => N663, Z => 
                           perm_output(158));
   C3536 : GTECH_XOR2 port map( A => plane1_2_60_port, B => N664, Z => 
                           perm_output(157));
   C3537 : GTECH_XOR2 port map( A => plane1_2_59_port, B => N665, Z => 
                           perm_output(156));
   C3538 : GTECH_XOR2 port map( A => plane1_2_58_port, B => N666, Z => 
                           perm_output(155));
   C3539 : GTECH_XOR2 port map( A => plane1_2_57_port, B => N667, Z => 
                           perm_output(154));
   C3540 : GTECH_XOR2 port map( A => plane1_2_56_port, B => N668, Z => 
                           perm_output(153));
   C3541 : GTECH_XOR2 port map( A => plane1_2_55_port, B => N669, Z => 
                           perm_output(152));
   C3542 : GTECH_XOR2 port map( A => plane1_2_54_port, B => N670, Z => 
                           perm_output(151));
   C3543 : GTECH_XOR2 port map( A => plane1_2_53_port, B => N671, Z => 
                           perm_output(150));
   C3544 : GTECH_XOR2 port map( A => plane1_2_52_port, B => N672, Z => 
                           perm_output(149));
   C3545 : GTECH_XOR2 port map( A => plane1_2_51_port, B => N673, Z => 
                           perm_output(148));
   C3546 : GTECH_XOR2 port map( A => plane1_2_50_port, B => N674, Z => 
                           perm_output(147));
   C3547 : GTECH_XOR2 port map( A => plane1_2_49_port, B => N675, Z => 
                           perm_output(146));
   C3548 : GTECH_XOR2 port map( A => plane1_2_48_port, B => N676, Z => 
                           perm_output(145));
   C3549 : GTECH_XOR2 port map( A => plane1_2_47_port, B => N677, Z => 
                           perm_output(144));
   C3550 : GTECH_XOR2 port map( A => plane1_2_46_port, B => N678, Z => 
                           perm_output(143));
   C3551 : GTECH_XOR2 port map( A => plane1_2_45_port, B => N679, Z => 
                           perm_output(142));
   C3552 : GTECH_XOR2 port map( A => plane1_2_44_port, B => N680, Z => 
                           perm_output(141));
   C3553 : GTECH_XOR2 port map( A => plane1_2_43_port, B => N681, Z => 
                           perm_output(140));
   C3554 : GTECH_XOR2 port map( A => plane1_2_42_port, B => N682, Z => 
                           perm_output(139));
   C3555 : GTECH_XOR2 port map( A => plane1_2_41_port, B => N683, Z => 
                           perm_output(138));
   C3556 : GTECH_XOR2 port map( A => plane1_2_40_port, B => N684, Z => 
                           perm_output(137));
   C3557 : GTECH_XOR2 port map( A => plane1_2_39_port, B => N685, Z => 
                           perm_output(136));
   C3558 : GTECH_XOR2 port map( A => plane1_2_38_port, B => N686, Z => 
                           perm_output(135));
   C3559 : GTECH_XOR2 port map( A => plane1_2_37_port, B => N687, Z => 
                           perm_output(134));
   C3560 : GTECH_XOR2 port map( A => plane1_2_36_port, B => N688, Z => 
                           perm_output(133));
   C3561 : GTECH_XOR2 port map( A => plane1_2_35_port, B => N689, Z => 
                           perm_output(132));
   C3562 : GTECH_XOR2 port map( A => plane1_2_34_port, B => N690, Z => 
                           perm_output(131));
   C3563 : GTECH_XOR2 port map( A => plane1_2_33_port, B => N691, Z => 
                           perm_output(130));
   C3564 : GTECH_XOR2 port map( A => plane1_2_32_port, B => N692, Z => 
                           perm_output(129));
   I_276 : GTECH_NOT port map( A => plane0_2_127_port, Z => N693);
   I_277 : GTECH_NOT port map( A => plane0_2_126_port, Z => N694);
   I_278 : GTECH_NOT port map( A => plane0_2_125_port, Z => N695);
   I_279 : GTECH_NOT port map( A => plane0_2_124_port, Z => N696);
   I_280 : GTECH_NOT port map( A => plane0_2_123_port, Z => N697);
   I_281 : GTECH_NOT port map( A => plane0_2_122_port, Z => N698);
   I_282 : GTECH_NOT port map( A => plane0_2_121_port, Z => N699);
   I_283 : GTECH_NOT port map( A => plane0_2_120_port, Z => N700);
   I_284 : GTECH_NOT port map( A => plane0_2_119_port, Z => N701);
   I_285 : GTECH_NOT port map( A => plane0_2_118_port, Z => N702);
   I_286 : GTECH_NOT port map( A => plane0_2_117_port, Z => N703);
   I_287 : GTECH_NOT port map( A => plane0_2_116_port, Z => N704);
   I_288 : GTECH_NOT port map( A => plane0_2_115_port, Z => N705);
   I_289 : GTECH_NOT port map( A => plane0_2_114_port, Z => N706);
   I_290 : GTECH_NOT port map( A => plane0_2_113_port, Z => N707);
   I_291 : GTECH_NOT port map( A => plane0_2_112_port, Z => N708);
   I_292 : GTECH_NOT port map( A => plane0_2_111_port, Z => N709);
   I_293 : GTECH_NOT port map( A => plane0_2_110_port, Z => N710);
   I_294 : GTECH_NOT port map( A => plane0_2_109_port, Z => N711);
   I_295 : GTECH_NOT port map( A => plane0_2_108_port, Z => N712);
   I_296 : GTECH_NOT port map( A => add_rnd_const_small_11_port, Z => N713);
   I_297 : GTECH_NOT port map( A => add_rnd_const_small_10_port, Z => N714);
   I_298 : GTECH_NOT port map( A => add_rnd_const_small_9_port, Z => N715);
   I_299 : GTECH_NOT port map( A => add_rnd_const_small_8_port, Z => N716);
   I_300 : GTECH_NOT port map( A => add_rnd_const_small_7_port, Z => N717);
   I_301 : GTECH_NOT port map( A => add_rnd_const_small_6_port, Z => N718);
   I_302 : GTECH_NOT port map( A => add_rnd_const_small_5_port, Z => N719);
   I_303 : GTECH_NOT port map( A => add_rnd_const_small_4_port, Z => N720);
   I_304 : GTECH_NOT port map( A => add_rnd_const_small_3_port, Z => N721);
   I_305 : GTECH_NOT port map( A => add_rnd_const_small_2_port, Z => N722);
   I_306 : GTECH_NOT port map( A => add_rnd_const_small_1_port, Z => N723);
   I_307 : GTECH_NOT port map( A => add_rnd_const_small_0_port, Z => N724);
   I_308 : GTECH_NOT port map( A => plane0_2_95_port, Z => N725);
   I_309 : GTECH_NOT port map( A => plane0_2_94_port, Z => N726);
   I_310 : GTECH_NOT port map( A => plane0_2_93_port, Z => N727);
   I_311 : GTECH_NOT port map( A => plane0_2_92_port, Z => N728);
   I_312 : GTECH_NOT port map( A => plane0_2_91_port, Z => N729);
   I_313 : GTECH_NOT port map( A => plane0_2_90_port, Z => N730);
   I_314 : GTECH_NOT port map( A => plane0_2_89_port, Z => N731);
   I_315 : GTECH_NOT port map( A => plane0_2_88_port, Z => N732);
   I_316 : GTECH_NOT port map( A => plane0_2_87_port, Z => N733);
   I_317 : GTECH_NOT port map( A => plane0_2_86_port, Z => N734);
   I_318 : GTECH_NOT port map( A => plane0_2_85_port, Z => N735);
   I_319 : GTECH_NOT port map( A => plane0_2_84_port, Z => N736);
   I_320 : GTECH_NOT port map( A => plane0_2_83_port, Z => N737);
   I_321 : GTECH_NOT port map( A => plane0_2_82_port, Z => N738);
   I_322 : GTECH_NOT port map( A => plane0_2_81_port, Z => N739);
   I_323 : GTECH_NOT port map( A => plane0_2_80_port, Z => N740);
   I_324 : GTECH_NOT port map( A => plane0_2_79_port, Z => N741);
   I_325 : GTECH_NOT port map( A => plane0_2_78_port, Z => N742);
   I_326 : GTECH_NOT port map( A => plane0_2_77_port, Z => N743);
   I_327 : GTECH_NOT port map( A => plane0_2_76_port, Z => N744);
   I_328 : GTECH_NOT port map( A => plane0_2_75_port, Z => N745);
   I_329 : GTECH_NOT port map( A => plane0_2_74_port, Z => N746);
   I_330 : GTECH_NOT port map( A => plane0_2_73_port, Z => N747);
   I_331 : GTECH_NOT port map( A => plane0_2_72_port, Z => N748);
   I_332 : GTECH_NOT port map( A => plane0_2_71_port, Z => N749);
   I_333 : GTECH_NOT port map( A => plane0_2_70_port, Z => N750);
   I_334 : GTECH_NOT port map( A => plane0_2_69_port, Z => N751);
   I_335 : GTECH_NOT port map( A => plane0_2_68_port, Z => N752);
   I_336 : GTECH_NOT port map( A => plane0_2_67_port, Z => N753);
   I_337 : GTECH_NOT port map( A => plane0_2_66_port, Z => N754);
   I_338 : GTECH_NOT port map( A => plane0_2_65_port, Z => N755);
   I_339 : GTECH_NOT port map( A => plane0_2_64_port, Z => N756);
   I_340 : GTECH_NOT port map( A => plane0_2_63_port, Z => N757);
   I_341 : GTECH_NOT port map( A => plane0_2_62_port, Z => N758);
   I_342 : GTECH_NOT port map( A => plane0_2_61_port, Z => N759);
   I_343 : GTECH_NOT port map( A => plane0_2_60_port, Z => N760);
   I_344 : GTECH_NOT port map( A => plane0_2_59_port, Z => N761);
   I_345 : GTECH_NOT port map( A => plane0_2_58_port, Z => N762);
   I_346 : GTECH_NOT port map( A => plane0_2_57_port, Z => N763);
   I_347 : GTECH_NOT port map( A => plane0_2_56_port, Z => N764);
   I_348 : GTECH_NOT port map( A => plane0_2_55_port, Z => N765);
   I_349 : GTECH_NOT port map( A => plane0_2_54_port, Z => N766);
   I_350 : GTECH_NOT port map( A => plane0_2_53_port, Z => N767);
   I_351 : GTECH_NOT port map( A => plane0_2_52_port, Z => N768);
   I_352 : GTECH_NOT port map( A => plane0_2_51_port, Z => N769);
   I_353 : GTECH_NOT port map( A => plane0_2_50_port, Z => N770);
   I_354 : GTECH_NOT port map( A => plane0_2_49_port, Z => N771);
   I_355 : GTECH_NOT port map( A => plane0_2_48_port, Z => N772);
   I_356 : GTECH_NOT port map( A => plane0_2_47_port, Z => N773);
   I_357 : GTECH_NOT port map( A => plane0_2_46_port, Z => N774);
   I_358 : GTECH_NOT port map( A => plane0_2_45_port, Z => N775);
   I_359 : GTECH_NOT port map( A => plane0_2_44_port, Z => N776);
   I_360 : GTECH_NOT port map( A => plane0_2_43_port, Z => N777);
   I_361 : GTECH_NOT port map( A => plane0_2_42_port, Z => N778);
   I_362 : GTECH_NOT port map( A => plane0_2_41_port, Z => N779);
   I_363 : GTECH_NOT port map( A => plane0_2_40_port, Z => N780);
   I_364 : GTECH_NOT port map( A => plane0_2_39_port, Z => N781);
   I_365 : GTECH_NOT port map( A => plane0_2_38_port, Z => N782);
   I_366 : GTECH_NOT port map( A => plane0_2_37_port, Z => N783);
   I_367 : GTECH_NOT port map( A => plane0_2_36_port, Z => N784);
   I_368 : GTECH_NOT port map( A => plane0_2_35_port, Z => N785);
   I_369 : GTECH_NOT port map( A => plane0_2_34_port, Z => N786);
   I_370 : GTECH_NOT port map( A => plane0_2_33_port, Z => N787);
   I_371 : GTECH_NOT port map( A => plane0_2_32_port, Z => N788);
   I_372 : GTECH_NOT port map( A => plane0_2_31_port, Z => N789);
   I_373 : GTECH_NOT port map( A => plane0_2_30_port, Z => N790);
   I_374 : GTECH_NOT port map( A => plane0_2_29_port, Z => N791);
   I_375 : GTECH_NOT port map( A => plane0_2_28_port, Z => N792);
   I_376 : GTECH_NOT port map( A => plane0_2_27_port, Z => N793);
   I_377 : GTECH_NOT port map( A => plane0_2_26_port, Z => N794);
   I_378 : GTECH_NOT port map( A => plane0_2_25_port, Z => N795);
   I_379 : GTECH_NOT port map( A => plane0_2_24_port, Z => N796);
   I_380 : GTECH_NOT port map( A => plane0_2_23_port, Z => N797);
   I_381 : GTECH_NOT port map( A => plane0_2_22_port, Z => N798);
   I_382 : GTECH_NOT port map( A => plane0_2_21_port, Z => N799);
   I_383 : GTECH_NOT port map( A => plane0_2_20_port, Z => N800);
   I_384 : GTECH_NOT port map( A => plane0_2_19_port, Z => N801);
   I_385 : GTECH_NOT port map( A => plane0_2_18_port, Z => N802);
   I_386 : GTECH_NOT port map( A => plane0_2_17_port, Z => N803);
   I_387 : GTECH_NOT port map( A => plane0_2_16_port, Z => N804);
   I_388 : GTECH_NOT port map( A => plane0_2_15_port, Z => N805);
   I_389 : GTECH_NOT port map( A => plane0_2_14_port, Z => N806);
   I_390 : GTECH_NOT port map( A => plane0_2_13_port, Z => N807);
   I_391 : GTECH_NOT port map( A => plane0_2_12_port, Z => N808);
   I_392 : GTECH_NOT port map( A => plane0_2_11_port, Z => N809);
   I_393 : GTECH_NOT port map( A => plane0_2_10_port, Z => N810);
   I_394 : GTECH_NOT port map( A => plane0_2_9_port, Z => N811);
   I_395 : GTECH_NOT port map( A => plane0_2_8_port, Z => N812);
   I_396 : GTECH_NOT port map( A => plane0_2_7_port, Z => N813);
   I_397 : GTECH_NOT port map( A => plane0_2_6_port, Z => N814);
   I_398 : GTECH_NOT port map( A => plane0_2_5_port, Z => N815);
   I_399 : GTECH_NOT port map( A => plane0_2_4_port, Z => N816);
   I_400 : GTECH_NOT port map( A => plane0_2_3_port, Z => N817);
   I_401 : GTECH_NOT port map( A => plane0_2_2_port, Z => N818);
   I_402 : GTECH_NOT port map( A => plane0_2_1_port, Z => N819);
   I_403 : GTECH_NOT port map( A => plane0_2_0_port, Z => N820);
   C3693 : GTECH_AND2 port map( A => N693, B => plane1_2_31_port, Z => N821);
   C3694 : GTECH_AND2 port map( A => N694, B => plane1_2_30_port, Z => N822);
   C3695 : GTECH_AND2 port map( A => N695, B => plane1_2_29_port, Z => N823);
   C3696 : GTECH_AND2 port map( A => N696, B => plane1_2_28_port, Z => N824);
   C3697 : GTECH_AND2 port map( A => N697, B => plane1_2_27_port, Z => N825);
   C3698 : GTECH_AND2 port map( A => N698, B => plane1_2_26_port, Z => N826);
   C3699 : GTECH_AND2 port map( A => N699, B => plane1_2_25_port, Z => N827);
   C3700 : GTECH_AND2 port map( A => N700, B => plane1_2_24_port, Z => N828);
   C3701 : GTECH_AND2 port map( A => N701, B => plane1_2_23_port, Z => N829);
   C3702 : GTECH_AND2 port map( A => N702, B => plane1_2_22_port, Z => N830);
   C3703 : GTECH_AND2 port map( A => N703, B => plane1_2_21_port, Z => N831);
   C3704 : GTECH_AND2 port map( A => N704, B => plane1_2_20_port, Z => N832);
   C3705 : GTECH_AND2 port map( A => N705, B => plane1_2_19_port, Z => N833);
   C3706 : GTECH_AND2 port map( A => N706, B => plane1_2_18_port, Z => N834);
   C3707 : GTECH_AND2 port map( A => N707, B => plane1_2_17_port, Z => N835);
   C3708 : GTECH_AND2 port map( A => N708, B => plane1_2_16_port, Z => N836);
   C3709 : GTECH_AND2 port map( A => N709, B => plane1_2_15_port, Z => N837);
   C3710 : GTECH_AND2 port map( A => N710, B => plane1_2_14_port, Z => N838);
   C3711 : GTECH_AND2 port map( A => N711, B => plane1_2_13_port, Z => N839);
   C3712 : GTECH_AND2 port map( A => N712, B => plane1_2_12_port, Z => N840);
   C3713 : GTECH_AND2 port map( A => N713, B => plane1_2_11_port, Z => N841);
   C3714 : GTECH_AND2 port map( A => N714, B => plane1_2_10_port, Z => N842);
   C3715 : GTECH_AND2 port map( A => N715, B => plane1_2_9_port, Z => N843);
   C3716 : GTECH_AND2 port map( A => N716, B => plane1_2_8_port, Z => N844);
   C3717 : GTECH_AND2 port map( A => N717, B => plane1_2_7_port, Z => N845);
   C3718 : GTECH_AND2 port map( A => N718, B => plane1_2_6_port, Z => N846);
   C3719 : GTECH_AND2 port map( A => N719, B => plane1_2_5_port, Z => N847);
   C3720 : GTECH_AND2 port map( A => N720, B => plane1_2_4_port, Z => N848);
   C3721 : GTECH_AND2 port map( A => N721, B => plane1_2_3_port, Z => N849);
   C3722 : GTECH_AND2 port map( A => N722, B => plane1_2_2_port, Z => N850);
   C3723 : GTECH_AND2 port map( A => N723, B => plane1_2_1_port, Z => N851);
   C3724 : GTECH_AND2 port map( A => N724, B => plane1_2_0_port, Z => N852);
   C3725 : GTECH_AND2 port map( A => N725, B => plane1_2_127_port, Z => N853);
   C3726 : GTECH_AND2 port map( A => N726, B => plane1_2_126_port, Z => N854);
   C3727 : GTECH_AND2 port map( A => N727, B => plane1_2_125_port, Z => N855);
   C3728 : GTECH_AND2 port map( A => N728, B => plane1_2_124_port, Z => N856);
   C3729 : GTECH_AND2 port map( A => N729, B => plane1_2_123_port, Z => N857);
   C3730 : GTECH_AND2 port map( A => N730, B => plane1_2_122_port, Z => N858);
   C3731 : GTECH_AND2 port map( A => N731, B => plane1_2_121_port, Z => N859);
   C3732 : GTECH_AND2 port map( A => N732, B => plane1_2_120_port, Z => N860);
   C3733 : GTECH_AND2 port map( A => N733, B => plane1_2_119_port, Z => N861);
   C3734 : GTECH_AND2 port map( A => N734, B => plane1_2_118_port, Z => N862);
   C3735 : GTECH_AND2 port map( A => N735, B => plane1_2_117_port, Z => N863);
   C3736 : GTECH_AND2 port map( A => N736, B => plane1_2_116_port, Z => N864);
   C3737 : GTECH_AND2 port map( A => N737, B => plane1_2_115_port, Z => N865);
   C3738 : GTECH_AND2 port map( A => N738, B => plane1_2_114_port, Z => N866);
   C3739 : GTECH_AND2 port map( A => N739, B => plane1_2_113_port, Z => N867);
   C3740 : GTECH_AND2 port map( A => N740, B => plane1_2_112_port, Z => N868);
   C3741 : GTECH_AND2 port map( A => N741, B => plane1_2_111_port, Z => N869);
   C3742 : GTECH_AND2 port map( A => N742, B => plane1_2_110_port, Z => N870);
   C3743 : GTECH_AND2 port map( A => N743, B => plane1_2_109_port, Z => N871);
   C3744 : GTECH_AND2 port map( A => N744, B => plane1_2_108_port, Z => N872);
   C3745 : GTECH_AND2 port map( A => N745, B => plane1_2_107_port, Z => N873);
   C3746 : GTECH_AND2 port map( A => N746, B => plane1_2_106_port, Z => N874);
   C3747 : GTECH_AND2 port map( A => N747, B => plane1_2_105_port, Z => N875);
   C3748 : GTECH_AND2 port map( A => N748, B => plane1_2_104_port, Z => N876);
   C3749 : GTECH_AND2 port map( A => N749, B => plane1_2_103_port, Z => N877);
   C3750 : GTECH_AND2 port map( A => N750, B => plane1_2_102_port, Z => N878);
   C3751 : GTECH_AND2 port map( A => N751, B => plane1_2_101_port, Z => N879);
   C3752 : GTECH_AND2 port map( A => N752, B => plane1_2_100_port, Z => N880);
   C3753 : GTECH_AND2 port map( A => N753, B => plane1_2_99_port, Z => N881);
   C3754 : GTECH_AND2 port map( A => N754, B => plane1_2_98_port, Z => N882);
   C3755 : GTECH_AND2 port map( A => N755, B => plane1_2_97_port, Z => N883);
   C3756 : GTECH_AND2 port map( A => N756, B => plane1_2_96_port, Z => N884);
   C3757 : GTECH_AND2 port map( A => N757, B => plane1_2_95_port, Z => N885);
   C3758 : GTECH_AND2 port map( A => N758, B => plane1_2_94_port, Z => N886);
   C3759 : GTECH_AND2 port map( A => N759, B => plane1_2_93_port, Z => N887);
   C3760 : GTECH_AND2 port map( A => N760, B => plane1_2_92_port, Z => N888);
   C3761 : GTECH_AND2 port map( A => N761, B => plane1_2_91_port, Z => N889);
   C3762 : GTECH_AND2 port map( A => N762, B => plane1_2_90_port, Z => N890);
   C3763 : GTECH_AND2 port map( A => N763, B => plane1_2_89_port, Z => N891);
   C3764 : GTECH_AND2 port map( A => N764, B => plane1_2_88_port, Z => N892);
   C3765 : GTECH_AND2 port map( A => N765, B => plane1_2_87_port, Z => N893);
   C3766 : GTECH_AND2 port map( A => N766, B => plane1_2_86_port, Z => N894);
   C3767 : GTECH_AND2 port map( A => N767, B => plane1_2_85_port, Z => N895);
   C3768 : GTECH_AND2 port map( A => N768, B => plane1_2_84_port, Z => N896);
   C3769 : GTECH_AND2 port map( A => N769, B => plane1_2_83_port, Z => N897);
   C3770 : GTECH_AND2 port map( A => N770, B => plane1_2_82_port, Z => N898);
   C3771 : GTECH_AND2 port map( A => N771, B => plane1_2_81_port, Z => N899);
   C3772 : GTECH_AND2 port map( A => N772, B => plane1_2_80_port, Z => N900);
   C3773 : GTECH_AND2 port map( A => N773, B => plane1_2_79_port, Z => N901);
   C3774 : GTECH_AND2 port map( A => N774, B => plane1_2_78_port, Z => N902);
   C3775 : GTECH_AND2 port map( A => N775, B => plane1_2_77_port, Z => N903);
   C3776 : GTECH_AND2 port map( A => N776, B => plane1_2_76_port, Z => N904);
   C3777 : GTECH_AND2 port map( A => N777, B => plane1_2_75_port, Z => N905);
   C3778 : GTECH_AND2 port map( A => N778, B => plane1_2_74_port, Z => N906);
   C3779 : GTECH_AND2 port map( A => N779, B => plane1_2_73_port, Z => N907);
   C3780 : GTECH_AND2 port map( A => N780, B => plane1_2_72_port, Z => N908);
   C3781 : GTECH_AND2 port map( A => N781, B => plane1_2_71_port, Z => N909);
   C3782 : GTECH_AND2 port map( A => N782, B => plane1_2_70_port, Z => N910);
   C3783 : GTECH_AND2 port map( A => N783, B => plane1_2_69_port, Z => N911);
   C3784 : GTECH_AND2 port map( A => N784, B => plane1_2_68_port, Z => N912);
   C3785 : GTECH_AND2 port map( A => N785, B => plane1_2_67_port, Z => N913);
   C3786 : GTECH_AND2 port map( A => N786, B => plane1_2_66_port, Z => N914);
   C3787 : GTECH_AND2 port map( A => N787, B => plane1_2_65_port, Z => N915);
   C3788 : GTECH_AND2 port map( A => N788, B => plane1_2_64_port, Z => N916);
   C3789 : GTECH_AND2 port map( A => N789, B => plane1_2_63_port, Z => N917);
   C3790 : GTECH_AND2 port map( A => N790, B => plane1_2_62_port, Z => N918);
   C3791 : GTECH_AND2 port map( A => N791, B => plane1_2_61_port, Z => N919);
   C3792 : GTECH_AND2 port map( A => N792, B => plane1_2_60_port, Z => N920);
   C3793 : GTECH_AND2 port map( A => N793, B => plane1_2_59_port, Z => N921);
   C3794 : GTECH_AND2 port map( A => N794, B => plane1_2_58_port, Z => N922);
   C3795 : GTECH_AND2 port map( A => N795, B => plane1_2_57_port, Z => N923);
   C3796 : GTECH_AND2 port map( A => N796, B => plane1_2_56_port, Z => N924);
   C3797 : GTECH_AND2 port map( A => N797, B => plane1_2_55_port, Z => N925);
   C3798 : GTECH_AND2 port map( A => N798, B => plane1_2_54_port, Z => N926);
   C3799 : GTECH_AND2 port map( A => N799, B => plane1_2_53_port, Z => N927);
   C3800 : GTECH_AND2 port map( A => N800, B => plane1_2_52_port, Z => N928);
   C3801 : GTECH_AND2 port map( A => N801, B => plane1_2_51_port, Z => N929);
   C3802 : GTECH_AND2 port map( A => N802, B => plane1_2_50_port, Z => N930);
   C3803 : GTECH_AND2 port map( A => N803, B => plane1_2_49_port, Z => N931);
   C3804 : GTECH_AND2 port map( A => N804, B => plane1_2_48_port, Z => N932);
   C3805 : GTECH_AND2 port map( A => N805, B => plane1_2_47_port, Z => N933);
   C3806 : GTECH_AND2 port map( A => N806, B => plane1_2_46_port, Z => N934);
   C3807 : GTECH_AND2 port map( A => N807, B => plane1_2_45_port, Z => N935);
   C3808 : GTECH_AND2 port map( A => N808, B => plane1_2_44_port, Z => N936);
   C3809 : GTECH_AND2 port map( A => N809, B => plane1_2_43_port, Z => N937);
   C3810 : GTECH_AND2 port map( A => N810, B => plane1_2_42_port, Z => N938);
   C3811 : GTECH_AND2 port map( A => N811, B => plane1_2_41_port, Z => N939);
   C3812 : GTECH_AND2 port map( A => N812, B => plane1_2_40_port, Z => N940);
   C3813 : GTECH_AND2 port map( A => N813, B => plane1_2_39_port, Z => N941);
   C3814 : GTECH_AND2 port map( A => N814, B => plane1_2_38_port, Z => N942);
   C3815 : GTECH_AND2 port map( A => N815, B => plane1_2_37_port, Z => N943);
   C3816 : GTECH_AND2 port map( A => N816, B => plane1_2_36_port, Z => N944);
   C3817 : GTECH_AND2 port map( A => N817, B => plane1_2_35_port, Z => N945);
   C3818 : GTECH_AND2 port map( A => N818, B => plane1_2_34_port, Z => N946);
   C3819 : GTECH_AND2 port map( A => N819, B => plane1_2_33_port, Z => N947);
   C3820 : GTECH_AND2 port map( A => N820, B => plane1_2_32_port, Z => N948);
   C3821 : GTECH_XOR2 port map( A => plane2_2_116_port, B => N821, Z => 
                           perm_output(295));
   C3822 : GTECH_XOR2 port map( A => plane2_2_115_port, B => N822, Z => 
                           perm_output(294));
   C3823 : GTECH_XOR2 port map( A => plane2_2_114_port, B => N823, Z => 
                           perm_output(293));
   C3824 : GTECH_XOR2 port map( A => plane2_2_113_port, B => N824, Z => 
                           perm_output(292));
   C3825 : GTECH_XOR2 port map( A => plane2_2_112_port, B => N825, Z => 
                           perm_output(291));
   C3826 : GTECH_XOR2 port map( A => plane2_2_111_port, B => N826, Z => 
                           perm_output(290));
   C3827 : GTECH_XOR2 port map( A => plane2_2_110_port, B => N827, Z => 
                           perm_output(289));
   C3828 : GTECH_XOR2 port map( A => plane2_2_109_port, B => N828, Z => 
                           perm_output(288));
   C3829 : GTECH_XOR2 port map( A => plane2_2_108_port, B => N829, Z => 
                           perm_output(319));
   C3830 : GTECH_XOR2 port map( A => plane2_2_107_port, B => N830, Z => 
                           perm_output(318));
   C3831 : GTECH_XOR2 port map( A => plane2_2_106_port, B => N831, Z => 
                           perm_output(317));
   C3832 : GTECH_XOR2 port map( A => plane2_2_105_port, B => N832, Z => 
                           perm_output(316));
   C3833 : GTECH_XOR2 port map( A => plane2_2_104_port, B => N833, Z => 
                           perm_output(315));
   C3834 : GTECH_XOR2 port map( A => plane2_2_103_port, B => N834, Z => 
                           perm_output(314));
   C3835 : GTECH_XOR2 port map( A => plane2_2_102_port, B => N835, Z => 
                           perm_output(313));
   C3836 : GTECH_XOR2 port map( A => plane2_2_101_port, B => N836, Z => 
                           perm_output(312));
   C3837 : GTECH_XOR2 port map( A => plane2_2_100_port, B => N837, Z => 
                           perm_output(311));
   C3838 : GTECH_XOR2 port map( A => plane2_2_99_port, B => N838, Z => 
                           perm_output(310));
   C3839 : GTECH_XOR2 port map( A => plane2_2_98_port, B => N839, Z => 
                           perm_output(309));
   C3840 : GTECH_XOR2 port map( A => plane2_2_97_port, B => N840, Z => 
                           perm_output(308));
   C3841 : GTECH_XOR2 port map( A => plane2_2_96_port, B => N841, Z => 
                           perm_output(307));
   C3842 : GTECH_XOR2 port map( A => plane2_2_127_port, B => N842, Z => 
                           perm_output(306));
   C3843 : GTECH_XOR2 port map( A => plane2_2_126_port, B => N843, Z => 
                           perm_output(305));
   C3844 : GTECH_XOR2 port map( A => plane2_2_125_port, B => N844, Z => 
                           perm_output(304));
   C3845 : GTECH_XOR2 port map( A => plane2_2_124_port, B => N845, Z => 
                           perm_output(303));
   C3846 : GTECH_XOR2 port map( A => plane2_2_123_port, B => N846, Z => 
                           perm_output(302));
   C3847 : GTECH_XOR2 port map( A => plane2_2_122_port, B => N847, Z => 
                           perm_output(301));
   C3848 : GTECH_XOR2 port map( A => plane2_2_121_port, B => N848, Z => 
                           perm_output(300));
   C3849 : GTECH_XOR2 port map( A => plane2_2_120_port, B => N849, Z => 
                           perm_output(299));
   C3850 : GTECH_XOR2 port map( A => plane2_2_119_port, B => N850, Z => 
                           perm_output(298));
   C3851 : GTECH_XOR2 port map( A => plane2_2_118_port, B => N851, Z => 
                           perm_output(297));
   C3852 : GTECH_XOR2 port map( A => plane2_2_117_port, B => N852, Z => 
                           perm_output(296));
   C3853 : GTECH_XOR2 port map( A => plane2_2_84_port, B => N853, Z => 
                           perm_output(263));
   C3854 : GTECH_XOR2 port map( A => plane2_2_83_port, B => N854, Z => 
                           perm_output(262));
   C3855 : GTECH_XOR2 port map( A => plane2_2_82_port, B => N855, Z => 
                           perm_output(261));
   C3856 : GTECH_XOR2 port map( A => plane2_2_81_port, B => N856, Z => 
                           perm_output(260));
   C3857 : GTECH_XOR2 port map( A => plane2_2_80_port, B => N857, Z => 
                           perm_output(259));
   C3858 : GTECH_XOR2 port map( A => plane2_2_79_port, B => N858, Z => 
                           perm_output(258));
   C3859 : GTECH_XOR2 port map( A => plane2_2_78_port, B => N859, Z => 
                           perm_output(257));
   C3860 : GTECH_XOR2 port map( A => plane2_2_77_port, B => N860, Z => 
                           perm_output(256));
   C3861 : GTECH_XOR2 port map( A => plane2_2_76_port, B => N861, Z => 
                           perm_output(287));
   C3862 : GTECH_XOR2 port map( A => plane2_2_75_port, B => N862, Z => 
                           perm_output(286));
   C3863 : GTECH_XOR2 port map( A => plane2_2_74_port, B => N863, Z => 
                           perm_output(285));
   C3864 : GTECH_XOR2 port map( A => plane2_2_73_port, B => N864, Z => 
                           perm_output(284));
   C3865 : GTECH_XOR2 port map( A => plane2_2_72_port, B => N865, Z => 
                           perm_output(283));
   C3866 : GTECH_XOR2 port map( A => plane2_2_71_port, B => N866, Z => 
                           perm_output(282));
   C3867 : GTECH_XOR2 port map( A => plane2_2_70_port, B => N867, Z => 
                           perm_output(281));
   C3868 : GTECH_XOR2 port map( A => plane2_2_69_port, B => N868, Z => 
                           perm_output(280));
   C3869 : GTECH_XOR2 port map( A => plane2_2_68_port, B => N869, Z => 
                           perm_output(279));
   C3870 : GTECH_XOR2 port map( A => plane2_2_67_port, B => N870, Z => 
                           perm_output(278));
   C3871 : GTECH_XOR2 port map( A => plane2_2_66_port, B => N871, Z => 
                           perm_output(277));
   C3872 : GTECH_XOR2 port map( A => plane2_2_65_port, B => N872, Z => 
                           perm_output(276));
   C3873 : GTECH_XOR2 port map( A => plane2_2_64_port, B => N873, Z => 
                           perm_output(275));
   C3874 : GTECH_XOR2 port map( A => plane2_2_95_port, B => N874, Z => 
                           perm_output(274));
   C3875 : GTECH_XOR2 port map( A => plane2_2_94_port, B => N875, Z => 
                           perm_output(273));
   C3876 : GTECH_XOR2 port map( A => plane2_2_93_port, B => N876, Z => 
                           perm_output(272));
   C3877 : GTECH_XOR2 port map( A => plane2_2_92_port, B => N877, Z => 
                           perm_output(271));
   C3878 : GTECH_XOR2 port map( A => plane2_2_91_port, B => N878, Z => 
                           perm_output(270));
   C3879 : GTECH_XOR2 port map( A => plane2_2_90_port, B => N879, Z => 
                           perm_output(269));
   C3880 : GTECH_XOR2 port map( A => plane2_2_89_port, B => N880, Z => 
                           perm_output(268));
   C3881 : GTECH_XOR2 port map( A => plane2_2_88_port, B => N881, Z => 
                           perm_output(267));
   C3882 : GTECH_XOR2 port map( A => plane2_2_87_port, B => N882, Z => 
                           perm_output(266));
   C3883 : GTECH_XOR2 port map( A => plane2_2_86_port, B => N883, Z => 
                           perm_output(265));
   C3884 : GTECH_XOR2 port map( A => plane2_2_85_port, B => N884, Z => 
                           perm_output(264));
   C3885 : GTECH_XOR2 port map( A => plane2_2_52_port, B => N885, Z => 
                           perm_output(359));
   C3886 : GTECH_XOR2 port map( A => plane2_2_51_port, B => N886, Z => 
                           perm_output(358));
   C3887 : GTECH_XOR2 port map( A => plane2_2_50_port, B => N887, Z => 
                           perm_output(357));
   C3888 : GTECH_XOR2 port map( A => plane2_2_49_port, B => N888, Z => 
                           perm_output(356));
   C3889 : GTECH_XOR2 port map( A => plane2_2_48_port, B => N889, Z => 
                           perm_output(355));
   C3890 : GTECH_XOR2 port map( A => plane2_2_47_port, B => N890, Z => 
                           perm_output(354));
   C3891 : GTECH_XOR2 port map( A => plane2_2_46_port, B => N891, Z => 
                           perm_output(353));
   C3892 : GTECH_XOR2 port map( A => plane2_2_45_port, B => N892, Z => 
                           perm_output(352));
   C3893 : GTECH_XOR2 port map( A => plane2_2_44_port, B => N893, Z => 
                           perm_output(383));
   C3894 : GTECH_XOR2 port map( A => plane2_2_43_port, B => N894, Z => 
                           perm_output(382));
   C3895 : GTECH_XOR2 port map( A => plane2_2_42_port, B => N895, Z => 
                           perm_output(381));
   C3896 : GTECH_XOR2 port map( A => plane2_2_41_port, B => N896, Z => 
                           perm_output(380));
   C3897 : GTECH_XOR2 port map( A => plane2_2_40_port, B => N897, Z => 
                           perm_output(379));
   C3898 : GTECH_XOR2 port map( A => plane2_2_39_port, B => N898, Z => 
                           perm_output(378));
   C3899 : GTECH_XOR2 port map( A => plane2_2_38_port, B => N899, Z => 
                           perm_output(377));
   C3900 : GTECH_XOR2 port map( A => plane2_2_37_port, B => N900, Z => 
                           perm_output(376));
   C3901 : GTECH_XOR2 port map( A => plane2_2_36_port, B => N901, Z => 
                           perm_output(375));
   C3902 : GTECH_XOR2 port map( A => plane2_2_35_port, B => N902, Z => 
                           perm_output(374));
   C3903 : GTECH_XOR2 port map( A => plane2_2_34_port, B => N903, Z => 
                           perm_output(373));
   C3904 : GTECH_XOR2 port map( A => plane2_2_33_port, B => N904, Z => 
                           perm_output(372));
   C3905 : GTECH_XOR2 port map( A => plane2_2_32_port, B => N905, Z => 
                           perm_output(371));
   C3906 : GTECH_XOR2 port map( A => plane2_2_63_port, B => N906, Z => 
                           perm_output(370));
   C3907 : GTECH_XOR2 port map( A => plane2_2_62_port, B => N907, Z => 
                           perm_output(369));
   C3908 : GTECH_XOR2 port map( A => plane2_2_61_port, B => N908, Z => 
                           perm_output(368));
   C3909 : GTECH_XOR2 port map( A => plane2_2_60_port, B => N909, Z => 
                           perm_output(367));
   C3910 : GTECH_XOR2 port map( A => plane2_2_59_port, B => N910, Z => 
                           perm_output(366));
   C3911 : GTECH_XOR2 port map( A => plane2_2_58_port, B => N911, Z => 
                           perm_output(365));
   C3912 : GTECH_XOR2 port map( A => plane2_2_57_port, B => N912, Z => 
                           perm_output(364));
   C3913 : GTECH_XOR2 port map( A => plane2_2_56_port, B => N913, Z => 
                           perm_output(363));
   C3914 : GTECH_XOR2 port map( A => plane2_2_55_port, B => N914, Z => 
                           perm_output(362));
   C3915 : GTECH_XOR2 port map( A => plane2_2_54_port, B => N915, Z => 
                           perm_output(361));
   C3916 : GTECH_XOR2 port map( A => plane2_2_53_port, B => N916, Z => 
                           perm_output(360));
   C3917 : GTECH_XOR2 port map( A => plane2_2_20_port, B => N917, Z => 
                           perm_output(327));
   C3918 : GTECH_XOR2 port map( A => plane2_2_19_port, B => N918, Z => 
                           perm_output(326));
   C3919 : GTECH_XOR2 port map( A => plane2_2_18_port, B => N919, Z => 
                           perm_output(325));
   C3920 : GTECH_XOR2 port map( A => plane2_2_17_port, B => N920, Z => 
                           perm_output(324));
   C3921 : GTECH_XOR2 port map( A => plane2_2_16_port, B => N921, Z => 
                           perm_output(323));
   C3922 : GTECH_XOR2 port map( A => plane2_2_15_port, B => N922, Z => 
                           perm_output(322));
   C3923 : GTECH_XOR2 port map( A => plane2_2_14_port, B => N923, Z => 
                           perm_output(321));
   C3924 : GTECH_XOR2 port map( A => plane2_2_13_port, B => N924, Z => 
                           perm_output(320));
   C3925 : GTECH_XOR2 port map( A => plane2_2_12_port, B => N925, Z => 
                           perm_output(351));
   C3926 : GTECH_XOR2 port map( A => plane2_2_11_port, B => N926, Z => 
                           perm_output(350));
   C3927 : GTECH_XOR2 port map( A => plane2_2_10_port, B => N927, Z => 
                           perm_output(349));
   C3928 : GTECH_XOR2 port map( A => plane2_2_9_port, B => N928, Z => 
                           perm_output(348));
   C3929 : GTECH_XOR2 port map( A => plane2_2_8_port, B => N929, Z => 
                           perm_output(347));
   C3930 : GTECH_XOR2 port map( A => plane2_2_7_port, B => N930, Z => 
                           perm_output(346));
   C3931 : GTECH_XOR2 port map( A => plane2_2_6_port, B => N931, Z => 
                           perm_output(345));
   C3932 : GTECH_XOR2 port map( A => plane2_2_5_port, B => N932, Z => 
                           perm_output(344));
   C3933 : GTECH_XOR2 port map( A => plane2_2_4_port, B => N933, Z => 
                           perm_output(343));
   C3934 : GTECH_XOR2 port map( A => plane2_2_3_port, B => N934, Z => 
                           perm_output(342));
   C3935 : GTECH_XOR2 port map( A => plane2_2_2_port, B => N935, Z => 
                           perm_output(341));
   C3936 : GTECH_XOR2 port map( A => plane2_2_1_port, B => N936, Z => 
                           perm_output(340));
   C3937 : GTECH_XOR2 port map( A => plane2_2_0_port, B => N937, Z => 
                           perm_output(339));
   C3938 : GTECH_XOR2 port map( A => plane2_2_31_port, B => N938, Z => 
                           perm_output(338));
   C3939 : GTECH_XOR2 port map( A => plane2_2_30_port, B => N939, Z => 
                           perm_output(337));
   C3940 : GTECH_XOR2 port map( A => plane2_2_29_port, B => N940, Z => 
                           perm_output(336));
   C3941 : GTECH_XOR2 port map( A => plane2_2_28_port, B => N941, Z => 
                           perm_output(335));
   C3942 : GTECH_XOR2 port map( A => plane2_2_27_port, B => N942, Z => 
                           perm_output(334));
   C3943 : GTECH_XOR2 port map( A => plane2_2_26_port, B => N943, Z => 
                           perm_output(333));
   C3944 : GTECH_XOR2 port map( A => plane2_2_25_port, B => N944, Z => 
                           perm_output(332));
   C3945 : GTECH_XOR2 port map( A => plane2_2_24_port, B => N945, Z => 
                           perm_output(331));
   C3946 : GTECH_XOR2 port map( A => plane2_2_23_port, B => N946, Z => 
                           perm_output(330));
   C3947 : GTECH_XOR2 port map( A => plane2_2_22_port, B => N947, Z => 
                           perm_output(329));
   C3948 : GTECH_XOR2 port map( A => plane2_2_21_port, B => N948, Z => 
                           perm_output(328));

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_LWC_1.all;

entity reg_custom_LEN128_1 is

   port( clk, en : in std_logic;  din : in std_logic_vector (127 downto 0);  
         qout : out std_logic_vector (127 downto 0));

end reg_custom_LEN128_1;

architecture SYN_RTL of reg_custom_LEN128_1 is
   
   component SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
      generic ( ac_as_q, ac_as_qn, sc_ss_q : integer );
      port(
         clear, preset, enable, data_in, synch_clear, synch_preset, 
            synch_toggle, synch_enable, next_state, clocked_on : in std_logic;
         Q, QN : buffer std_logic
      );
   end component;
   
   signal X_Logic0_port, clk_port, en_port, din_127_port, din_126_port, 
      din_125_port, din_124_port, din_123_port, din_122_port, din_121_port, 
      din_120_port, din_119_port, din_118_port, din_117_port, din_116_port, 
      din_115_port, din_114_port, din_113_port, din_112_port, din_111_port, 
      din_110_port, din_109_port, din_108_port, din_107_port, din_106_port, 
      din_105_port, din_104_port, din_103_port, din_102_port, din_101_port, 
      din_100_port, din_99_port, din_98_port, din_97_port, din_96_port, 
      din_95_port, din_94_port, din_93_port, din_92_port, din_91_port, 
      din_90_port, din_89_port, din_88_port, din_87_port, din_86_port, 
      din_85_port, din_84_port, din_83_port, din_82_port, din_81_port, 
      din_80_port, din_79_port, din_78_port, din_77_port, din_76_port, 
      din_75_port, din_74_port, din_73_port, din_72_port, din_71_port, 
      din_70_port, din_69_port, din_68_port, din_67_port, din_66_port, 
      din_65_port, din_64_port, din_63_port, din_62_port, din_61_port, 
      din_60_port, din_59_port, din_58_port, din_57_port, din_56_port, 
      din_55_port, din_54_port, din_53_port, din_52_port, din_51_port, 
      din_50_port, din_49_port, din_48_port, din_47_port, din_46_port, 
      din_45_port, din_44_port, din_43_port, din_42_port, din_41_port, 
      din_40_port, din_39_port, din_38_port, din_37_port, din_36_port, 
      din_35_port, din_34_port, din_33_port, din_32_port, din_31_port, 
      din_30_port, din_29_port, din_28_port, din_27_port, din_26_port, 
      din_25_port, din_24_port, din_23_port, din_22_port, din_21_port, 
      din_20_port, din_19_port, din_18_port, din_17_port, din_16_port, 
      din_15_port, din_14_port, din_13_port, din_12_port, din_11_port, 
      din_10_port, din_9_port, din_8_port, din_7_port, din_6_port, din_5_port, 
      din_4_port, din_3_port, din_2_port, din_1_port, din_0_port, qout_127_port
      , qout_126_port, qout_125_port, qout_124_port, qout_123_port, 
      qout_122_port, qout_121_port, qout_120_port, qout_119_port, qout_118_port
      , qout_117_port, qout_116_port, qout_115_port, qout_114_port, 
      qout_113_port, qout_112_port, qout_111_port, qout_110_port, qout_109_port
      , qout_108_port, qout_107_port, qout_106_port, qout_105_port, 
      qout_104_port, qout_103_port, qout_102_port, qout_101_port, qout_100_port
      , qout_99_port, qout_98_port, qout_97_port, qout_96_port, qout_95_port, 
      qout_94_port, qout_93_port, qout_92_port, qout_91_port, qout_90_port, 
      qout_89_port, qout_88_port, qout_87_port, qout_86_port, qout_85_port, 
      qout_84_port, qout_83_port, qout_82_port, qout_81_port, qout_80_port, 
      qout_79_port, qout_78_port, qout_77_port, qout_76_port, qout_75_port, 
      qout_74_port, qout_73_port, qout_72_port, qout_71_port, qout_70_port, 
      qout_69_port, qout_68_port, qout_67_port, qout_66_port, qout_65_port, 
      qout_64_port, qout_63_port, qout_62_port, qout_61_port, qout_60_port, 
      qout_59_port, qout_58_port, qout_57_port, qout_56_port, qout_55_port, 
      qout_54_port, qout_53_port, qout_52_port, qout_51_port, qout_50_port, 
      qout_49_port, qout_48_port, qout_47_port, qout_46_port, qout_45_port, 
      qout_44_port, qout_43_port, qout_42_port, qout_41_port, qout_40_port, 
      qout_39_port, qout_38_port, qout_37_port, qout_36_port, qout_35_port, 
      qout_34_port, qout_33_port, qout_32_port, qout_31_port, qout_30_port, 
      qout_29_port, qout_28_port, qout_27_port, qout_26_port, qout_25_port, 
      qout_24_port, qout_23_port, qout_22_port, qout_21_port, qout_20_port, 
      qout_19_port, qout_18_port, qout_17_port, qout_16_port, qout_15_port, 
      qout_14_port, qout_13_port, qout_12_port, qout_11_port, qout_10_port, 
      qout_9_port, qout_8_port, qout_7_port, qout_6_port, qout_5_port, 
      qout_4_port, qout_3_port, qout_2_port, qout_1_port, qout_0_port, n_1000, 
      n_1001, n_1002, n_1003, n_1004, n_1005, n_1006, n_1007, n_1008, n_1009, 
      n_1010, n_1011, n_1012, n_1013, n_1014, n_1015, n_1016, n_1017, n_1018, 
      n_1019, n_1020, n_1021, n_1022, n_1023, n_1024, n_1025, n_1026, n_1027, 
      n_1028, n_1029, n_1030, n_1031, n_1032, n_1033, n_1034, n_1035, n_1036, 
      n_1037, n_1038, n_1039, n_1040, n_1041, n_1042, n_1043, n_1044, n_1045, 
      n_1046, n_1047, n_1048, n_1049, n_1050, n_1051, n_1052, n_1053, n_1054, 
      n_1055, n_1056, n_1057, n_1058, n_1059, n_1060, n_1061, n_1062, n_1063, 
      n_1064, n_1065, n_1066, n_1067, n_1068, n_1069, n_1070, n_1071, n_1072, 
      n_1073, n_1074, n_1075, n_1076, n_1077, n_1078, n_1079, n_1080, n_1081, 
      n_1082, n_1083, n_1084, n_1085, n_1086, n_1087, n_1088, n_1089, n_1090, 
      n_1091, n_1092, n_1093, n_1094, n_1095, n_1096, n_1097, n_1098, n_1099, 
      n_1100, n_1101, n_1102, n_1103, n_1104, n_1105, n_1106, n_1107, n_1108, 
      n_1109, n_1110, n_1111, n_1112, n_1113, n_1114, n_1115, n_1116, n_1117, 
      n_1118, n_1119, n_1120, n_1121, n_1122, n_1123, n_1124, n_1125, n_1126, 
      n_1127 : std_logic;

begin
   clk_port <= clk;
   en_port <= en;
   ( din_127_port, din_126_port, din_125_port, din_124_port, din_123_port, 
      din_122_port, din_121_port, din_120_port, din_119_port, din_118_port, 
      din_117_port, din_116_port, din_115_port, din_114_port, din_113_port, 
      din_112_port, din_111_port, din_110_port, din_109_port, din_108_port, 
      din_107_port, din_106_port, din_105_port, din_104_port, din_103_port, 
      din_102_port, din_101_port, din_100_port, din_99_port, din_98_port, 
      din_97_port, din_96_port, din_95_port, din_94_port, din_93_port, 
      din_92_port, din_91_port, din_90_port, din_89_port, din_88_port, 
      din_87_port, din_86_port, din_85_port, din_84_port, din_83_port, 
      din_82_port, din_81_port, din_80_port, din_79_port, din_78_port, 
      din_77_port, din_76_port, din_75_port, din_74_port, din_73_port, 
      din_72_port, din_71_port, din_70_port, din_69_port, din_68_port, 
      din_67_port, din_66_port, din_65_port, din_64_port, din_63_port, 
      din_62_port, din_61_port, din_60_port, din_59_port, din_58_port, 
      din_57_port, din_56_port, din_55_port, din_54_port, din_53_port, 
      din_52_port, din_51_port, din_50_port, din_49_port, din_48_port, 
      din_47_port, din_46_port, din_45_port, din_44_port, din_43_port, 
      din_42_port, din_41_port, din_40_port, din_39_port, din_38_port, 
      din_37_port, din_36_port, din_35_port, din_34_port, din_33_port, 
      din_32_port, din_31_port, din_30_port, din_29_port, din_28_port, 
      din_27_port, din_26_port, din_25_port, din_24_port, din_23_port, 
      din_22_port, din_21_port, din_20_port, din_19_port, din_18_port, 
      din_17_port, din_16_port, din_15_port, din_14_port, din_13_port, 
      din_12_port, din_11_port, din_10_port, din_9_port, din_8_port, din_7_port
      , din_6_port, din_5_port, din_4_port, din_3_port, din_2_port, din_1_port,
      din_0_port ) <= din;
   qout <= ( qout_127_port, qout_126_port, qout_125_port, qout_124_port, 
      qout_123_port, qout_122_port, qout_121_port, qout_120_port, qout_119_port
      , qout_118_port, qout_117_port, qout_116_port, qout_115_port, 
      qout_114_port, qout_113_port, qout_112_port, qout_111_port, qout_110_port
      , qout_109_port, qout_108_port, qout_107_port, qout_106_port, 
      qout_105_port, qout_104_port, qout_103_port, qout_102_port, qout_101_port
      , qout_100_port, qout_99_port, qout_98_port, qout_97_port, qout_96_port, 
      qout_95_port, qout_94_port, qout_93_port, qout_92_port, qout_91_port, 
      qout_90_port, qout_89_port, qout_88_port, qout_87_port, qout_86_port, 
      qout_85_port, qout_84_port, qout_83_port, qout_82_port, qout_81_port, 
      qout_80_port, qout_79_port, qout_78_port, qout_77_port, qout_76_port, 
      qout_75_port, qout_74_port, qout_73_port, qout_72_port, qout_71_port, 
      qout_70_port, qout_69_port, qout_68_port, qout_67_port, qout_66_port, 
      qout_65_port, qout_64_port, qout_63_port, qout_62_port, qout_61_port, 
      qout_60_port, qout_59_port, qout_58_port, qout_57_port, qout_56_port, 
      qout_55_port, qout_54_port, qout_53_port, qout_52_port, qout_51_port, 
      qout_50_port, qout_49_port, qout_48_port, qout_47_port, qout_46_port, 
      qout_45_port, qout_44_port, qout_43_port, qout_42_port, qout_41_port, 
      qout_40_port, qout_39_port, qout_38_port, qout_37_port, qout_36_port, 
      qout_35_port, qout_34_port, qout_33_port, qout_32_port, qout_31_port, 
      qout_30_port, qout_29_port, qout_28_port, qout_27_port, qout_26_port, 
      qout_25_port, qout_24_port, qout_23_port, qout_22_port, qout_21_port, 
      qout_20_port, qout_19_port, qout_18_port, qout_17_port, qout_16_port, 
      qout_15_port, qout_14_port, qout_13_port, qout_12_port, qout_11_port, 
      qout_10_port, qout_9_port, qout_8_port, qout_7_port, qout_6_port, 
      qout_5_port, qout_4_port, qout_3_port, qout_2_port, qout_1_port, 
      qout_0_port );
   
   qout_reg_127_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_127_port, clocked_on => clk_port, Q => qout_127_port, QN => 
               n_1000);
   qout_reg_126_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_126_port, clocked_on => clk_port, Q => qout_126_port, QN => 
               n_1001);
   qout_reg_125_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_125_port, clocked_on => clk_port, Q => qout_125_port, QN => 
               n_1002);
   qout_reg_124_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_124_port, clocked_on => clk_port, Q => qout_124_port, QN => 
               n_1003);
   qout_reg_123_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_123_port, clocked_on => clk_port, Q => qout_123_port, QN => 
               n_1004);
   qout_reg_122_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_122_port, clocked_on => clk_port, Q => qout_122_port, QN => 
               n_1005);
   qout_reg_121_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_121_port, clocked_on => clk_port, Q => qout_121_port, QN => 
               n_1006);
   qout_reg_120_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_120_port, clocked_on => clk_port, Q => qout_120_port, QN => 
               n_1007);
   qout_reg_119_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_119_port, clocked_on => clk_port, Q => qout_119_port, QN => 
               n_1008);
   qout_reg_118_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_118_port, clocked_on => clk_port, Q => qout_118_port, QN => 
               n_1009);
   qout_reg_117_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_117_port, clocked_on => clk_port, Q => qout_117_port, QN => 
               n_1010);
   qout_reg_116_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_116_port, clocked_on => clk_port, Q => qout_116_port, QN => 
               n_1011);
   qout_reg_115_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_115_port, clocked_on => clk_port, Q => qout_115_port, QN => 
               n_1012);
   qout_reg_114_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_114_port, clocked_on => clk_port, Q => qout_114_port, QN => 
               n_1013);
   qout_reg_113_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_113_port, clocked_on => clk_port, Q => qout_113_port, QN => 
               n_1014);
   qout_reg_112_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_112_port, clocked_on => clk_port, Q => qout_112_port, QN => 
               n_1015);
   qout_reg_111_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_111_port, clocked_on => clk_port, Q => qout_111_port, QN => 
               n_1016);
   qout_reg_110_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_110_port, clocked_on => clk_port, Q => qout_110_port, QN => 
               n_1017);
   qout_reg_109_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_109_port, clocked_on => clk_port, Q => qout_109_port, QN => 
               n_1018);
   qout_reg_108_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_108_port, clocked_on => clk_port, Q => qout_108_port, QN => 
               n_1019);
   qout_reg_107_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_107_port, clocked_on => clk_port, Q => qout_107_port, QN => 
               n_1020);
   qout_reg_106_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_106_port, clocked_on => clk_port, Q => qout_106_port, QN => 
               n_1021);
   qout_reg_105_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_105_port, clocked_on => clk_port, Q => qout_105_port, QN => 
               n_1022);
   qout_reg_104_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_104_port, clocked_on => clk_port, Q => qout_104_port, QN => 
               n_1023);
   qout_reg_103_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_103_port, clocked_on => clk_port, Q => qout_103_port, QN => 
               n_1024);
   qout_reg_102_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_102_port, clocked_on => clk_port, Q => qout_102_port, QN => 
               n_1025);
   qout_reg_101_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_101_port, clocked_on => clk_port, Q => qout_101_port, QN => 
               n_1026);
   qout_reg_100_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_100_port, clocked_on => clk_port, Q => qout_100_port, QN => 
               n_1027);
   qout_reg_99_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_99_port, clocked_on => clk_port, Q => qout_99_port, QN => 
               n_1028);
   qout_reg_98_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_98_port, clocked_on => clk_port, Q => qout_98_port, QN => 
               n_1029);
   qout_reg_97_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_97_port, clocked_on => clk_port, Q => qout_97_port, QN => 
               n_1030);
   qout_reg_96_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_96_port, clocked_on => clk_port, Q => qout_96_port, QN => 
               n_1031);
   qout_reg_95_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_95_port, clocked_on => clk_port, Q => qout_95_port, QN => 
               n_1032);
   qout_reg_94_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_94_port, clocked_on => clk_port, Q => qout_94_port, QN => 
               n_1033);
   qout_reg_93_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_93_port, clocked_on => clk_port, Q => qout_93_port, QN => 
               n_1034);
   qout_reg_92_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_92_port, clocked_on => clk_port, Q => qout_92_port, QN => 
               n_1035);
   qout_reg_91_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_91_port, clocked_on => clk_port, Q => qout_91_port, QN => 
               n_1036);
   qout_reg_90_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_90_port, clocked_on => clk_port, Q => qout_90_port, QN => 
               n_1037);
   qout_reg_89_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_89_port, clocked_on => clk_port, Q => qout_89_port, QN => 
               n_1038);
   qout_reg_88_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_88_port, clocked_on => clk_port, Q => qout_88_port, QN => 
               n_1039);
   qout_reg_87_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_87_port, clocked_on => clk_port, Q => qout_87_port, QN => 
               n_1040);
   qout_reg_86_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_86_port, clocked_on => clk_port, Q => qout_86_port, QN => 
               n_1041);
   qout_reg_85_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_85_port, clocked_on => clk_port, Q => qout_85_port, QN => 
               n_1042);
   qout_reg_84_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_84_port, clocked_on => clk_port, Q => qout_84_port, QN => 
               n_1043);
   qout_reg_83_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_83_port, clocked_on => clk_port, Q => qout_83_port, QN => 
               n_1044);
   qout_reg_82_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_82_port, clocked_on => clk_port, Q => qout_82_port, QN => 
               n_1045);
   qout_reg_81_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_81_port, clocked_on => clk_port, Q => qout_81_port, QN => 
               n_1046);
   qout_reg_80_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_80_port, clocked_on => clk_port, Q => qout_80_port, QN => 
               n_1047);
   qout_reg_79_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_79_port, clocked_on => clk_port, Q => qout_79_port, QN => 
               n_1048);
   qout_reg_78_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_78_port, clocked_on => clk_port, Q => qout_78_port, QN => 
               n_1049);
   qout_reg_77_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_77_port, clocked_on => clk_port, Q => qout_77_port, QN => 
               n_1050);
   qout_reg_76_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_76_port, clocked_on => clk_port, Q => qout_76_port, QN => 
               n_1051);
   qout_reg_75_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_75_port, clocked_on => clk_port, Q => qout_75_port, QN => 
               n_1052);
   qout_reg_74_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_74_port, clocked_on => clk_port, Q => qout_74_port, QN => 
               n_1053);
   qout_reg_73_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_73_port, clocked_on => clk_port, Q => qout_73_port, QN => 
               n_1054);
   qout_reg_72_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_72_port, clocked_on => clk_port, Q => qout_72_port, QN => 
               n_1055);
   qout_reg_71_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_71_port, clocked_on => clk_port, Q => qout_71_port, QN => 
               n_1056);
   qout_reg_70_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_70_port, clocked_on => clk_port, Q => qout_70_port, QN => 
               n_1057);
   qout_reg_69_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_69_port, clocked_on => clk_port, Q => qout_69_port, QN => 
               n_1058);
   qout_reg_68_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_68_port, clocked_on => clk_port, Q => qout_68_port, QN => 
               n_1059);
   qout_reg_67_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_67_port, clocked_on => clk_port, Q => qout_67_port, QN => 
               n_1060);
   qout_reg_66_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_66_port, clocked_on => clk_port, Q => qout_66_port, QN => 
               n_1061);
   qout_reg_65_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_65_port, clocked_on => clk_port, Q => qout_65_port, QN => 
               n_1062);
   qout_reg_64_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_64_port, clocked_on => clk_port, Q => qout_64_port, QN => 
               n_1063);
   qout_reg_63_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_63_port, clocked_on => clk_port, Q => qout_63_port, QN => 
               n_1064);
   qout_reg_62_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_62_port, clocked_on => clk_port, Q => qout_62_port, QN => 
               n_1065);
   qout_reg_61_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_61_port, clocked_on => clk_port, Q => qout_61_port, QN => 
               n_1066);
   qout_reg_60_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_60_port, clocked_on => clk_port, Q => qout_60_port, QN => 
               n_1067);
   qout_reg_59_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_59_port, clocked_on => clk_port, Q => qout_59_port, QN => 
               n_1068);
   qout_reg_58_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_58_port, clocked_on => clk_port, Q => qout_58_port, QN => 
               n_1069);
   qout_reg_57_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_57_port, clocked_on => clk_port, Q => qout_57_port, QN => 
               n_1070);
   qout_reg_56_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_56_port, clocked_on => clk_port, Q => qout_56_port, QN => 
               n_1071);
   qout_reg_55_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_55_port, clocked_on => clk_port, Q => qout_55_port, QN => 
               n_1072);
   qout_reg_54_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_54_port, clocked_on => clk_port, Q => qout_54_port, QN => 
               n_1073);
   qout_reg_53_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_53_port, clocked_on => clk_port, Q => qout_53_port, QN => 
               n_1074);
   qout_reg_52_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_52_port, clocked_on => clk_port, Q => qout_52_port, QN => 
               n_1075);
   qout_reg_51_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_51_port, clocked_on => clk_port, Q => qout_51_port, QN => 
               n_1076);
   qout_reg_50_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_50_port, clocked_on => clk_port, Q => qout_50_port, QN => 
               n_1077);
   qout_reg_49_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_49_port, clocked_on => clk_port, Q => qout_49_port, QN => 
               n_1078);
   qout_reg_48_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_48_port, clocked_on => clk_port, Q => qout_48_port, QN => 
               n_1079);
   qout_reg_47_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_47_port, clocked_on => clk_port, Q => qout_47_port, QN => 
               n_1080);
   qout_reg_46_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_46_port, clocked_on => clk_port, Q => qout_46_port, QN => 
               n_1081);
   qout_reg_45_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_45_port, clocked_on => clk_port, Q => qout_45_port, QN => 
               n_1082);
   qout_reg_44_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_44_port, clocked_on => clk_port, Q => qout_44_port, QN => 
               n_1083);
   qout_reg_43_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_43_port, clocked_on => clk_port, Q => qout_43_port, QN => 
               n_1084);
   qout_reg_42_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_42_port, clocked_on => clk_port, Q => qout_42_port, QN => 
               n_1085);
   qout_reg_41_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_41_port, clocked_on => clk_port, Q => qout_41_port, QN => 
               n_1086);
   qout_reg_40_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_40_port, clocked_on => clk_port, Q => qout_40_port, QN => 
               n_1087);
   qout_reg_39_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_39_port, clocked_on => clk_port, Q => qout_39_port, QN => 
               n_1088);
   qout_reg_38_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_38_port, clocked_on => clk_port, Q => qout_38_port, QN => 
               n_1089);
   qout_reg_37_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_37_port, clocked_on => clk_port, Q => qout_37_port, QN => 
               n_1090);
   qout_reg_36_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_36_port, clocked_on => clk_port, Q => qout_36_port, QN => 
               n_1091);
   qout_reg_35_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_35_port, clocked_on => clk_port, Q => qout_35_port, QN => 
               n_1092);
   qout_reg_34_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_34_port, clocked_on => clk_port, Q => qout_34_port, QN => 
               n_1093);
   qout_reg_33_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_33_port, clocked_on => clk_port, Q => qout_33_port, QN => 
               n_1094);
   qout_reg_32_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_32_port, clocked_on => clk_port, Q => qout_32_port, QN => 
               n_1095);
   qout_reg_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_31_port, clocked_on => clk_port, Q => qout_31_port, QN => 
               n_1096);
   qout_reg_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_30_port, clocked_on => clk_port, Q => qout_30_port, QN => 
               n_1097);
   qout_reg_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_29_port, clocked_on => clk_port, Q => qout_29_port, QN => 
               n_1098);
   qout_reg_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_28_port, clocked_on => clk_port, Q => qout_28_port, QN => 
               n_1099);
   qout_reg_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_27_port, clocked_on => clk_port, Q => qout_27_port, QN => 
               n_1100);
   qout_reg_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_26_port, clocked_on => clk_port, Q => qout_26_port, QN => 
               n_1101);
   qout_reg_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_25_port, clocked_on => clk_port, Q => qout_25_port, QN => 
               n_1102);
   qout_reg_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_24_port, clocked_on => clk_port, Q => qout_24_port, QN => 
               n_1103);
   qout_reg_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_23_port, clocked_on => clk_port, Q => qout_23_port, QN => 
               n_1104);
   qout_reg_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_22_port, clocked_on => clk_port, Q => qout_22_port, QN => 
               n_1105);
   qout_reg_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_21_port, clocked_on => clk_port, Q => qout_21_port, QN => 
               n_1106);
   qout_reg_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_20_port, clocked_on => clk_port, Q => qout_20_port, QN => 
               n_1107);
   qout_reg_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_19_port, clocked_on => clk_port, Q => qout_19_port, QN => 
               n_1108);
   qout_reg_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_18_port, clocked_on => clk_port, Q => qout_18_port, QN => 
               n_1109);
   qout_reg_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_17_port, clocked_on => clk_port, Q => qout_17_port, QN => 
               n_1110);
   qout_reg_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_16_port, clocked_on => clk_port, Q => qout_16_port, QN => 
               n_1111);
   qout_reg_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_15_port, clocked_on => clk_port, Q => qout_15_port, QN => 
               n_1112);
   qout_reg_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_14_port, clocked_on => clk_port, Q => qout_14_port, QN => 
               n_1113);
   qout_reg_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_13_port, clocked_on => clk_port, Q => qout_13_port, QN => 
               n_1114);
   qout_reg_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_12_port, clocked_on => clk_port, Q => qout_12_port, QN => 
               n_1115);
   qout_reg_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_11_port, clocked_on => clk_port, Q => qout_11_port, QN => 
               n_1116);
   qout_reg_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => 
               din_10_port, clocked_on => clk_port, Q => qout_10_port, QN => 
               n_1117);
   qout_reg_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => din_9_port
               , clocked_on => clk_port, Q => qout_9_port, QN => n_1118);
   qout_reg_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => din_8_port
               , clocked_on => clk_port, Q => qout_8_port, QN => n_1119);
   qout_reg_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => din_7_port
               , clocked_on => clk_port, Q => qout_7_port, QN => n_1120);
   qout_reg_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => din_6_port
               , clocked_on => clk_port, Q => qout_6_port, QN => n_1121);
   qout_reg_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => din_5_port
               , clocked_on => clk_port, Q => qout_5_port, QN => n_1122);
   qout_reg_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => din_4_port
               , clocked_on => clk_port, Q => qout_4_port, QN => n_1123);
   qout_reg_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => din_3_port
               , clocked_on => clk_port, Q => qout_3_port, QN => n_1124);
   qout_reg_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => din_2_port
               , clocked_on => clk_port, Q => qout_2_port, QN => n_1125);
   qout_reg_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => din_1_port
               , clocked_on => clk_port, Q => qout_1_port, QN => n_1126);
   qout_reg_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => en_port, next_state => din_0_port
               , clocked_on => clk_port, Q => qout_0_port, QN => n_1127);
   X_Logic0_port <= '0';

end SYN_RTL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_LWC_1.all;

entity DATA_SIPO_2 is

   port( clk, rst, end_of_input : in std_logic;  data_p : out std_logic_vector 
         (31 downto 0);  data_valid_p : out std_logic;  data_ready_p : in 
         std_logic;  data_s : in std_logic_vector (31 downto 0);  data_valid_s 
         : in std_logic;  data_ready_s : out std_logic);

end DATA_SIPO_2;

architecture SYN_behavioral of DATA_SIPO_2 is

begin
   data_p <= ( data_s(31), data_s(30), data_s(29), data_s(28), data_s(27), 
      data_s(26), data_s(25), data_s(24), data_s(23), data_s(22), data_s(21), 
      data_s(20), data_s(19), data_s(18), data_s(17), data_s(16), data_s(15), 
      data_s(14), data_s(13), data_s(12), data_s(11), data_s(10), data_s(9), 
      data_s(8), data_s(7), data_s(6), data_s(5), data_s(4), data_s(3), 
      data_s(2), data_s(1), data_s(0) );
   data_valid_p <= data_valid_s;
   data_ready_s <= data_ready_p;

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_LWC_1.all;

entity cyclist_ops_DATA_LEN32_1 is

   port( clk, key_en : in std_logic;  state_main_en : in std_logic_vector (2 
         downto 0);  state_main_sel : in std_logic_vector (6 downto 0);  
         cyc_state_update_sel, xor_sel : in std_logic;  cycd_sel : in 
         std_logic_vector (1 downto 0);  extract_sel : in std_logic;  bdi_key :
         in std_logic_vector (31 downto 0);  cu_cd : in std_logic_vector (7 
         downto 0);  dcount_in, rnd_counter : in std_logic_vector (3 downto 0);
         bdo_out : out std_logic_vector (31 downto 0));

end cyclist_ops_DATA_LEN32_1;

architecture SYN_Behavioral of cyclist_ops_DATA_LEN32_1 is

   component GTECH_NOT
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component GTECH_XOR2
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component GTECH_BUF
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component xoodoo_round_ADDRESS_LEN384_1
      port( INPUT : in std_logic_vector (383 downto 0);  perm_output : out 
            std_logic_vector (383 downto 0);  RNDCTR : in std_logic_vector (3 
            downto 0));
   end component;
   
   component reg_custom_LEN128_1
      port( clk, en : in std_logic;  din : in std_logic_vector (127 downto 0); 
            qout : out std_logic_vector (127 downto 0));
   end component;
   
   component GTECH_AND2
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component GTECH_OR2
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15,
      N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30
      , N31, X_Logic1_port, X_Logic0_port, bdi_key_31_port, bdi_key_30_port, 
      bdi_key_29_port, bdi_key_28_port, bdi_key_27_port, bdi_key_26_port, 
      bdi_key_25_port, bdi_key_24_port, bdi_key_23_port, bdi_key_22_port, 
      bdi_key_21_port, bdi_key_20_port, bdi_key_19_port, bdi_key_18_port, 
      bdi_key_17_port, bdi_key_16_port, bdi_key_15_port, bdi_key_14_port, 
      bdi_key_13_port, bdi_key_12_port, bdi_key_11_port, bdi_key_10_port, 
      bdi_key_9_port, bdi_key_8_port, bdi_key_7_port, bdi_key_6_port, 
      bdi_key_5_port, bdi_key_4_port, bdi_key_3_port, bdi_key_2_port, 
      bdi_key_1_port, bdi_key_0_port, bdo_out_31_port, bdo_out_30_port, 
      bdo_out_29_port, bdo_out_28_port, bdo_out_27_port, bdo_out_26_port, 
      bdo_out_25_port, bdo_out_24_port, bdo_out_23_port, bdo_out_22_port, 
      bdo_out_21_port, bdo_out_20_port, bdo_out_19_port, bdo_out_18_port, 
      bdo_out_17_port, bdo_out_16_port, bdo_out_15_port, bdo_out_14_port, 
      bdo_out_13_port, bdo_out_12_port, bdo_out_11_port, bdo_out_10_port, 
      bdo_out_9_port, bdo_out_8_port, bdo_out_7_port, bdo_out_6_port, 
      bdo_out_5_port, bdo_out_4_port, bdo_out_3_port, bdo_out_2_port, 
      bdo_out_1_port, bdo_out_0_port, N32, N33, plane_x_127_port, 
      plane_x_126_port, plane_x_125_port, plane_x_124_port, plane_x_123_port, 
      plane_x_122_port, plane_x_121_port, plane_x_120_port, plane_x_119_port, 
      plane_x_118_port, plane_x_117_port, plane_x_116_port, plane_x_115_port, 
      plane_x_114_port, plane_x_113_port, plane_x_112_port, plane_x_111_port, 
      plane_x_110_port, plane_x_109_port, plane_x_108_port, plane_x_107_port, 
      plane_x_106_port, plane_x_105_port, plane_x_104_port, plane_x_103_port, 
      plane_x_102_port, plane_x_101_port, plane_x_100_port, plane_x_99_port, 
      plane_x_98_port, plane_x_97_port, plane_x_96_port, plane_x_95_port, 
      plane_x_94_port, plane_x_93_port, plane_x_92_port, plane_x_91_port, 
      plane_x_90_port, plane_x_89_port, plane_x_88_port, plane_x_87_port, 
      plane_x_86_port, plane_x_85_port, plane_x_84_port, plane_x_83_port, 
      plane_x_82_port, plane_x_81_port, plane_x_80_port, plane_x_79_port, 
      plane_x_78_port, plane_x_77_port, plane_x_76_port, plane_x_75_port, 
      plane_x_74_port, plane_x_73_port, plane_x_72_port, plane_x_71_port, 
      plane_x_70_port, plane_x_69_port, plane_x_68_port, plane_x_67_port, 
      plane_x_66_port, plane_x_65_port, plane_x_64_port, plane_x_63_port, 
      plane_x_62_port, plane_x_61_port, plane_x_60_port, plane_x_59_port, 
      plane_x_58_port, plane_x_57_port, plane_x_56_port, plane_x_55_port, 
      plane_x_54_port, plane_x_53_port, plane_x_52_port, plane_x_51_port, 
      plane_x_50_port, plane_x_49_port, plane_x_48_port, plane_x_47_port, 
      plane_x_46_port, plane_x_45_port, plane_x_44_port, plane_x_43_port, 
      plane_x_42_port, plane_x_41_port, plane_x_40_port, plane_x_39_port, 
      plane_x_38_port, plane_x_37_port, plane_x_36_port, plane_x_35_port, 
      plane_x_34_port, plane_x_33_port, plane_x_32_port, plane_x_31_port, 
      plane_x_30_port, plane_x_29_port, plane_x_28_port, plane_x_27_port, 
      plane_x_26_port, plane_x_25_port, plane_x_24_port, plane_x_23_port, 
      plane_x_22_port, plane_x_21_port, plane_x_20_port, plane_x_19_port, 
      plane_x_18_port, plane_x_17_port, plane_x_16_port, plane_x_15_port, 
      plane_x_14_port, plane_x_13_port, plane_x_12_port, plane_x_11_port, 
      plane_x_10_port, plane_x_9_port, plane_x_8_port, plane_x_7_port, 
      plane_x_6_port, plane_x_5_port, plane_x_4_port, plane_x_3_port, 
      plane_x_2_port, plane_x_1_port, plane_x_0_port, 
      state_main_out_plane0_127_port, state_main_out_plane0_126_port, 
      state_main_out_plane0_125_port, state_main_out_plane0_124_port, 
      state_main_out_plane0_123_port, state_main_out_plane0_122_port, 
      state_main_out_plane0_121_port, state_main_out_plane0_120_port, 
      state_main_out_plane0_119_port, state_main_out_plane0_118_port, 
      state_main_out_plane0_117_port, state_main_out_plane0_116_port, 
      state_main_out_plane0_115_port, state_main_out_plane0_114_port, 
      state_main_out_plane0_113_port, state_main_out_plane0_112_port, 
      state_main_out_plane0_111_port, state_main_out_plane0_110_port, 
      state_main_out_plane0_109_port, state_main_out_plane0_108_port, 
      state_main_out_plane0_107_port, state_main_out_plane0_106_port, 
      state_main_out_plane0_105_port, state_main_out_plane0_104_port, 
      state_main_out_plane0_103_port, state_main_out_plane0_102_port, 
      state_main_out_plane0_101_port, state_main_out_plane0_100_port, 
      state_main_out_plane0_99_port, state_main_out_plane0_98_port, 
      state_main_out_plane0_97_port, state_main_out_plane0_96_port, 
      state_main_out_plane0_95_port, state_main_out_plane0_94_port, 
      state_main_out_plane0_93_port, state_main_out_plane0_92_port, 
      state_main_out_plane0_91_port, state_main_out_plane0_90_port, 
      state_main_out_plane0_89_port, state_main_out_plane0_88_port, 
      state_main_out_plane0_87_port, state_main_out_plane0_86_port, 
      state_main_out_plane0_85_port, state_main_out_plane0_84_port, 
      state_main_out_plane0_83_port, state_main_out_plane0_82_port, 
      state_main_out_plane0_81_port, state_main_out_plane0_80_port, 
      state_main_out_plane0_79_port, state_main_out_plane0_78_port, 
      state_main_out_plane0_77_port, state_main_out_plane0_76_port, 
      state_main_out_plane0_75_port, state_main_out_plane0_74_port, 
      state_main_out_plane0_73_port, state_main_out_plane0_72_port, 
      state_main_out_plane0_71_port, state_main_out_plane0_70_port, 
      state_main_out_plane0_69_port, state_main_out_plane0_68_port, 
      state_main_out_plane0_67_port, state_main_out_plane0_66_port, 
      state_main_out_plane0_65_port, state_main_out_plane0_64_port, 
      state_main_out_plane0_63_port, state_main_out_plane0_62_port, 
      state_main_out_plane0_61_port, state_main_out_plane0_60_port, 
      state_main_out_plane0_59_port, state_main_out_plane0_58_port, 
      state_main_out_plane0_57_port, state_main_out_plane0_56_port, 
      state_main_out_plane0_55_port, state_main_out_plane0_54_port, 
      state_main_out_plane0_53_port, state_main_out_plane0_52_port, 
      state_main_out_plane0_51_port, state_main_out_plane0_50_port, 
      state_main_out_plane0_49_port, state_main_out_plane0_48_port, 
      state_main_out_plane0_47_port, state_main_out_plane0_46_port, 
      state_main_out_plane0_45_port, state_main_out_plane0_44_port, 
      state_main_out_plane0_43_port, state_main_out_plane0_42_port, 
      state_main_out_plane0_41_port, state_main_out_plane0_40_port, 
      state_main_out_plane0_39_port, state_main_out_plane0_38_port, 
      state_main_out_plane0_37_port, state_main_out_plane0_36_port, 
      state_main_out_plane0_35_port, state_main_out_plane0_34_port, 
      state_main_out_plane0_33_port, state_main_out_plane0_32_port, 
      state_main_out_plane0_31_port, state_main_out_plane0_30_port, 
      state_main_out_plane0_29_port, state_main_out_plane0_28_port, 
      state_main_out_plane0_27_port, state_main_out_plane0_26_port, 
      state_main_out_plane0_25_port, state_main_out_plane0_24_port, 
      state_main_out_plane0_23_port, state_main_out_plane0_22_port, 
      state_main_out_plane0_21_port, state_main_out_plane0_20_port, 
      state_main_out_plane0_19_port, state_main_out_plane0_18_port, 
      state_main_out_plane0_17_port, state_main_out_plane0_16_port, 
      state_main_out_plane0_15_port, state_main_out_plane0_14_port, 
      state_main_out_plane0_13_port, state_main_out_plane0_12_port, 
      state_main_out_plane0_11_port, state_main_out_plane0_10_port, 
      state_main_out_plane0_9_port, state_main_out_plane0_8_port, 
      state_main_out_plane0_7_port, state_main_out_plane0_6_port, 
      state_main_out_plane0_5_port, state_main_out_plane0_4_port, 
      state_main_out_plane0_3_port, state_main_out_plane0_2_port, 
      state_main_out_plane0_1_port, state_main_out_plane0_0_port, 
      state_main_out_plane1_127_port, state_main_out_plane1_126_port, 
      state_main_out_plane1_125_port, state_main_out_plane1_124_port, 
      state_main_out_plane1_123_port, state_main_out_plane1_122_port, 
      state_main_out_plane1_121_port, state_main_out_plane1_120_port, 
      state_main_out_plane1_119_port, state_main_out_plane1_118_port, 
      state_main_out_plane1_117_port, state_main_out_plane1_116_port, 
      state_main_out_plane1_115_port, state_main_out_plane1_114_port, 
      state_main_out_plane1_113_port, state_main_out_plane1_112_port, 
      state_main_out_plane1_111_port, state_main_out_plane1_110_port, 
      state_main_out_plane1_109_port, state_main_out_plane1_108_port, 
      state_main_out_plane1_107_port, state_main_out_plane1_106_port, 
      state_main_out_plane1_105_port, state_main_out_plane1_104_port, 
      state_main_out_plane1_103_port, state_main_out_plane1_102_port, 
      state_main_out_plane1_101_port, state_main_out_plane1_100_port, 
      state_main_out_plane1_99_port, state_main_out_plane1_98_port, 
      state_main_out_plane1_97_port, state_main_out_plane1_96_port, 
      state_main_out_plane1_95_port, state_main_out_plane1_94_port, 
      state_main_out_plane1_93_port, state_main_out_plane1_92_port, 
      state_main_out_plane1_91_port, state_main_out_plane1_90_port, 
      state_main_out_plane1_89_port, state_main_out_plane1_88_port, 
      state_main_out_plane1_87_port, state_main_out_plane1_86_port, 
      state_main_out_plane1_85_port, state_main_out_plane1_84_port, 
      state_main_out_plane1_83_port, state_main_out_plane1_82_port, 
      state_main_out_plane1_81_port, state_main_out_plane1_80_port, 
      state_main_out_plane1_79_port, state_main_out_plane1_78_port, 
      state_main_out_plane1_77_port, state_main_out_plane1_76_port, 
      state_main_out_plane1_75_port, state_main_out_plane1_74_port, 
      state_main_out_plane1_73_port, state_main_out_plane1_72_port, 
      state_main_out_plane1_71_port, state_main_out_plane1_70_port, 
      state_main_out_plane1_69_port, state_main_out_plane1_68_port, 
      state_main_out_plane1_67_port, state_main_out_plane1_66_port, 
      state_main_out_plane1_65_port, state_main_out_plane1_64_port, 
      state_main_out_plane1_63_port, state_main_out_plane1_62_port, 
      state_main_out_plane1_61_port, state_main_out_plane1_60_port, 
      state_main_out_plane1_59_port, state_main_out_plane1_58_port, 
      state_main_out_plane1_57_port, state_main_out_plane1_56_port, 
      state_main_out_plane1_55_port, state_main_out_plane1_54_port, 
      state_main_out_plane1_53_port, state_main_out_plane1_52_port, 
      state_main_out_plane1_51_port, state_main_out_plane1_50_port, 
      state_main_out_plane1_49_port, state_main_out_plane1_48_port, 
      state_main_out_plane1_47_port, state_main_out_plane1_46_port, 
      state_main_out_plane1_45_port, state_main_out_plane1_44_port, 
      state_main_out_plane1_43_port, state_main_out_plane1_42_port, 
      state_main_out_plane1_41_port, state_main_out_plane1_40_port, 
      state_main_out_plane1_39_port, state_main_out_plane1_38_port, 
      state_main_out_plane1_37_port, state_main_out_plane1_36_port, 
      state_main_out_plane1_35_port, state_main_out_plane1_34_port, 
      state_main_out_plane1_33_port, state_main_out_plane1_32_port, 
      state_main_out_plane1_31_port, state_main_out_plane1_30_port, 
      state_main_out_plane1_29_port, state_main_out_plane1_28_port, 
      state_main_out_plane1_27_port, state_main_out_plane1_26_port, 
      state_main_out_plane1_25_port, state_main_out_plane1_24_port, 
      state_main_out_plane1_23_port, state_main_out_plane1_22_port, 
      state_main_out_plane1_21_port, state_main_out_plane1_20_port, 
      state_main_out_plane1_19_port, state_main_out_plane1_18_port, 
      state_main_out_plane1_17_port, state_main_out_plane1_16_port, 
      state_main_out_plane1_15_port, state_main_out_plane1_14_port, 
      state_main_out_plane1_13_port, state_main_out_plane1_12_port, 
      state_main_out_plane1_11_port, state_main_out_plane1_10_port, 
      state_main_out_plane1_9_port, state_main_out_plane1_8_port, 
      state_main_out_plane1_7_port, state_main_out_plane1_6_port, 
      state_main_out_plane1_5_port, state_main_out_plane1_4_port, 
      state_main_out_plane1_3_port, state_main_out_plane1_2_port, 
      state_main_out_plane1_1_port, state_main_out_plane1_0_port, N34, N35, N36
      , N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, 
      N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65
      , N66, N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78, N79, 
      N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91, N92, N93, N94
      , N95, N96, N97, N98, N99, N100, N101, N102, N103, N104, N105, N106, N107
      , N108, N109, N110, N111, N112, N113, N114, N115, N116, N117, N118, N119,
      N120, N121, N122, N123, N124, N125, N126, N127, N128, N129, N130, N131, 
      N132, N133, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143, 
      N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154, N155, 
      N156, N157, N158, N159, N160, N161, state_main_out_plane2_127_port, 
      state_main_out_plane2_126_port, state_main_out_plane2_125_port, 
      state_main_out_plane2_124_port, state_main_out_plane2_123_port, 
      state_main_out_plane2_122_port, state_main_out_plane2_121_port, 
      state_main_out_plane2_120_port, state_main_out_plane2_119_port, 
      state_main_out_plane2_118_port, state_main_out_plane2_117_port, 
      state_main_out_plane2_116_port, state_main_out_plane2_115_port, 
      state_main_out_plane2_114_port, state_main_out_plane2_113_port, 
      state_main_out_plane2_112_port, state_main_out_plane2_111_port, 
      state_main_out_plane2_110_port, state_main_out_plane2_109_port, 
      state_main_out_plane2_108_port, state_main_out_plane2_107_port, 
      state_main_out_plane2_106_port, state_main_out_plane2_105_port, 
      state_main_out_plane2_104_port, state_main_out_plane2_103_port, 
      state_main_out_plane2_102_port, state_main_out_plane2_101_port, 
      state_main_out_plane2_100_port, state_main_out_plane2_99_port, 
      state_main_out_plane2_98_port, state_main_out_plane2_97_port, 
      state_main_out_plane2_96_port, state_main_out_plane2_95_port, 
      state_main_out_plane2_94_port, state_main_out_plane2_93_port, 
      state_main_out_plane2_92_port, state_main_out_plane2_91_port, 
      state_main_out_plane2_90_port, state_main_out_plane2_89_port, 
      state_main_out_plane2_88_port, state_main_out_plane2_87_port, 
      state_main_out_plane2_86_port, state_main_out_plane2_85_port, 
      state_main_out_plane2_84_port, state_main_out_plane2_83_port, 
      state_main_out_plane2_82_port, state_main_out_plane2_81_port, 
      state_main_out_plane2_80_port, state_main_out_plane2_79_port, 
      state_main_out_plane2_78_port, state_main_out_plane2_77_port, 
      state_main_out_plane2_76_port, state_main_out_plane2_75_port, 
      state_main_out_plane2_74_port, state_main_out_plane2_73_port, 
      state_main_out_plane2_72_port, state_main_out_plane2_71_port, 
      state_main_out_plane2_70_port, state_main_out_plane2_69_port, 
      state_main_out_plane2_68_port, state_main_out_plane2_67_port, 
      state_main_out_plane2_66_port, state_main_out_plane2_65_port, 
      state_main_out_plane2_64_port, state_main_out_plane2_63_port, 
      state_main_out_plane2_62_port, state_main_out_plane2_61_port, 
      state_main_out_plane2_60_port, state_main_out_plane2_59_port, 
      state_main_out_plane2_58_port, state_main_out_plane2_57_port, 
      state_main_out_plane2_56_port, state_main_out_plane2_55_port, 
      state_main_out_plane2_54_port, state_main_out_plane2_53_port, 
      state_main_out_plane2_52_port, state_main_out_plane2_51_port, 
      state_main_out_plane2_50_port, state_main_out_plane2_49_port, 
      state_main_out_plane2_48_port, state_main_out_plane2_47_port, 
      state_main_out_plane2_46_port, state_main_out_plane2_45_port, 
      state_main_out_plane2_44_port, state_main_out_plane2_43_port, 
      state_main_out_plane2_42_port, state_main_out_plane2_41_port, 
      state_main_out_plane2_40_port, state_main_out_plane2_39_port, 
      state_main_out_plane2_38_port, state_main_out_plane2_37_port, 
      state_main_out_plane2_36_port, state_main_out_plane2_35_port, 
      state_main_out_plane2_34_port, state_main_out_plane2_33_port, 
      state_main_out_plane2_32_port, state_main_out_plane2_31_port, 
      state_main_out_plane2_30_port, state_main_out_plane2_29_port, 
      state_main_out_plane2_28_port, state_main_out_plane2_27_port, 
      state_main_out_plane2_26_port, state_main_out_plane2_25_port, 
      state_main_out_plane2_24_port, state_main_out_plane2_23_port, 
      state_main_out_plane2_22_port, state_main_out_plane2_21_port, 
      state_main_out_plane2_20_port, state_main_out_plane2_19_port, 
      state_main_out_plane2_18_port, state_main_out_plane2_17_port, 
      state_main_out_plane2_16_port, state_main_out_plane2_15_port, 
      state_main_out_plane2_14_port, state_main_out_plane2_13_port, 
      state_main_out_plane2_12_port, state_main_out_plane2_11_port, 
      state_main_out_plane2_10_port, state_main_out_plane2_9_port, 
      state_main_out_plane2_8_port, state_main_out_plane2_7_port, 
      state_main_out_plane2_6_port, state_main_out_plane2_5_port, 
      state_main_out_plane2_4_port, state_main_out_plane2_3_port, 
      state_main_out_plane2_2_port, state_main_out_plane2_1_port, 
      state_main_out_plane2_0_port, N162, N163, N164, N165, N166, N167, N168, 
      N169, cycd_add_24_port, cycd_add_23_port, cycd_add_22_port, 
      cycd_add_21_port, cycd_add_20_port, cycd_add_19_port, cycd_add_18_port, 
      cycd_add_17_port, cycd_add_16_port, cycd_add_15_port, cycd_add_14_port, 
      cycd_add_13_port, cycd_add_12_port, cycd_add_11_port, cycd_add_10_port, 
      cycd_add_9_port, cycd_add_8_port, cycd_add_7_port, cycd_add_6_port, 
      cycd_add_5_port, cycd_add_4_port, cycd_add_3_port, cycd_add_2_port, 
      cycd_add_1_port, cycd_add_0_port, xor_mux_o_31_port, xor_mux_o_30_port, 
      xor_mux_o_29_port, xor_mux_o_28_port, xor_mux_o_27_port, 
      xor_mux_o_26_port, xor_mux_o_25_port, xor_mux_o_24_port, 
      xor_mux_o_23_port, xor_mux_o_22_port, xor_mux_o_21_port, 
      xor_mux_o_20_port, xor_mux_o_19_port, xor_mux_o_18_port, 
      xor_mux_o_17_port, xor_mux_o_16_port, xor_mux_o_15_port, 
      xor_mux_o_14_port, xor_mux_o_13_port, xor_mux_o_12_port, 
      xor_mux_o_11_port, xor_mux_o_10_port, xor_mux_o_9_port, xor_mux_o_8_port,
      xor_mux_o_7_port, xor_mux_o_6_port, xor_mux_o_5_port, xor_mux_o_4_port, 
      xor_mux_o_3_port, xor_mux_o_2_port, xor_mux_o_1_port, xor_mux_o_0_port, 
      temp_ram_31_port, temp_ram_30_port, temp_ram_29_port, temp_ram_28_port, 
      temp_ram_27_port, temp_ram_26_port, temp_ram_25_port, temp_ram_24_port, 
      temp_ram_23_port, temp_ram_22_port, temp_ram_21_port, temp_ram_20_port, 
      temp_ram_19_port, temp_ram_18_port, temp_ram_17_port, temp_ram_16_port, 
      temp_ram_15_port, temp_ram_14_port, temp_ram_13_port, temp_ram_12_port, 
      temp_ram_11_port, temp_ram_10_port, temp_ram_9_port, temp_ram_8_port, 
      temp_ram_7_port, temp_ram_6_port, temp_ram_5_port, temp_ram_4_port, 
      temp_ram_3_port, temp_ram_2_port, temp_ram_1_port, temp_ram_0_port, 
      temp_xor_out_31_port, temp_xor_out_30_port, temp_xor_out_29_port, 
      temp_xor_out_28_port, temp_xor_out_27_port, temp_xor_out_26_port, 
      temp_xor_out_25_port, temp_xor_out_24_port, temp_xor_out_23_port, 
      temp_xor_out_22_port, temp_xor_out_21_port, temp_xor_out_20_port, 
      temp_xor_out_19_port, temp_xor_out_18_port, temp_xor_out_17_port, 
      temp_xor_out_16_port, temp_xor_out_15_port, temp_xor_out_14_port, 
      temp_xor_out_13_port, temp_xor_out_12_port, temp_xor_out_11_port, 
      temp_xor_out_10_port, temp_xor_out_9_port, temp_xor_out_8_port, 
      temp_xor_out_7_port, temp_xor_out_6_port, temp_xor_out_5_port, 
      temp_xor_out_4_port, temp_xor_out_3_port, temp_xor_out_2_port, 
      temp_xor_out_1_port, temp_xor_out_0_port, N170, N171, N172, N173, N174, 
      N175, N176, N177, N178, decrypt_mux_31_port, decrypt_mux_30_port, 
      decrypt_mux_29_port, decrypt_mux_28_port, decrypt_mux_27_port, 
      decrypt_mux_26_port, decrypt_mux_25_port, decrypt_mux_24_port, 
      decrypt_mux_23_port, decrypt_mux_22_port, decrypt_mux_21_port, 
      decrypt_mux_20_port, decrypt_mux_19_port, decrypt_mux_18_port, 
      decrypt_mux_17_port, decrypt_mux_16_port, decrypt_mux_15_port, 
      decrypt_mux_14_port, decrypt_mux_13_port, decrypt_mux_12_port, 
      decrypt_mux_11_port, decrypt_mux_10_port, decrypt_mux_9_port, 
      decrypt_mux_8_port, N179, N180, temp_cyc_state_31_port, 
      temp_cyc_state_30_port, temp_cyc_state_29_port, temp_cyc_state_28_port, 
      temp_cyc_state_27_port, temp_cyc_state_26_port, temp_cyc_state_25_port, 
      temp_cyc_state_24_port, temp_cyc_state_23_port, temp_cyc_state_22_port, 
      temp_cyc_state_21_port, temp_cyc_state_20_port, temp_cyc_state_19_port, 
      temp_cyc_state_18_port, temp_cyc_state_17_port, temp_cyc_state_16_port, 
      temp_cyc_state_15_port, temp_cyc_state_14_port, temp_cyc_state_13_port, 
      temp_cyc_state_12_port, temp_cyc_state_11_port, temp_cyc_state_10_port, 
      temp_cyc_state_9_port, temp_cyc_state_8_port, temp_cyc_state_7_port, 
      temp_cyc_state_6_port, temp_cyc_state_5_port, temp_cyc_state_4_port, 
      temp_cyc_state_3_port, temp_cyc_state_2_port, temp_cyc_state_1_port, 
      temp_cyc_state_0_port, cyc_state_update_127_port, 
      cyc_state_update_126_port, cyc_state_update_125_port, 
      cyc_state_update_124_port, cyc_state_update_123_port, 
      cyc_state_update_122_port, cyc_state_update_121_port, 
      cyc_state_update_120_port, cyc_state_update_119_port, 
      cyc_state_update_118_port, cyc_state_update_117_port, 
      cyc_state_update_116_port, cyc_state_update_115_port, 
      cyc_state_update_114_port, cyc_state_update_113_port, 
      cyc_state_update_112_port, cyc_state_update_111_port, 
      cyc_state_update_110_port, cyc_state_update_109_port, 
      cyc_state_update_108_port, cyc_state_update_107_port, 
      cyc_state_update_106_port, cyc_state_update_105_port, 
      cyc_state_update_104_port, cyc_state_update_103_port, 
      cyc_state_update_102_port, cyc_state_update_101_port, 
      cyc_state_update_100_port, cyc_state_update_99_port, 
      cyc_state_update_98_port, cyc_state_update_97_port, 
      cyc_state_update_96_port, cyc_state_update_95_port, 
      cyc_state_update_94_port, cyc_state_update_93_port, 
      cyc_state_update_92_port, cyc_state_update_91_port, 
      cyc_state_update_90_port, cyc_state_update_89_port, 
      cyc_state_update_88_port, cyc_state_update_87_port, 
      cyc_state_update_86_port, cyc_state_update_85_port, 
      cyc_state_update_84_port, cyc_state_update_83_port, 
      cyc_state_update_82_port, cyc_state_update_81_port, 
      cyc_state_update_80_port, cyc_state_update_79_port, 
      cyc_state_update_78_port, cyc_state_update_77_port, 
      cyc_state_update_76_port, cyc_state_update_75_port, 
      cyc_state_update_74_port, cyc_state_update_73_port, 
      cyc_state_update_72_port, cyc_state_update_71_port, 
      cyc_state_update_70_port, cyc_state_update_69_port, 
      cyc_state_update_68_port, cyc_state_update_67_port, 
      cyc_state_update_66_port, cyc_state_update_65_port, 
      cyc_state_update_64_port, cyc_state_update_63_port, 
      cyc_state_update_62_port, cyc_state_update_61_port, 
      cyc_state_update_60_port, cyc_state_update_59_port, 
      cyc_state_update_58_port, cyc_state_update_57_port, 
      cyc_state_update_56_port, cyc_state_update_55_port, 
      cyc_state_update_54_port, cyc_state_update_53_port, 
      cyc_state_update_52_port, cyc_state_update_51_port, 
      cyc_state_update_50_port, cyc_state_update_49_port, 
      cyc_state_update_48_port, cyc_state_update_47_port, 
      cyc_state_update_46_port, cyc_state_update_45_port, 
      cyc_state_update_44_port, cyc_state_update_43_port, 
      cyc_state_update_42_port, cyc_state_update_41_port, 
      cyc_state_update_40_port, cyc_state_update_39_port, 
      cyc_state_update_38_port, cyc_state_update_37_port, 
      cyc_state_update_36_port, cyc_state_update_35_port, 
      cyc_state_update_34_port, cyc_state_update_33_port, 
      cyc_state_update_32_port, cyc_state_update_31_port, 
      cyc_state_update_30_port, cyc_state_update_29_port, 
      cyc_state_update_28_port, cyc_state_update_27_port, 
      cyc_state_update_26_port, cyc_state_update_25_port, 
      cyc_state_update_24_port, cyc_state_update_23_port, 
      cyc_state_update_22_port, cyc_state_update_21_port, 
      cyc_state_update_20_port, cyc_state_update_19_port, 
      cyc_state_update_18_port, cyc_state_update_17_port, 
      cyc_state_update_16_port, cyc_state_update_15_port, 
      cyc_state_update_14_port, cyc_state_update_13_port, 
      cyc_state_update_12_port, cyc_state_update_11_port, 
      cyc_state_update_10_port, cyc_state_update_9_port, 
      cyc_state_update_8_port, cyc_state_update_7_port, cyc_state_update_6_port
      , cyc_state_update_5_port, cyc_state_update_4_port, 
      cyc_state_update_3_port, cyc_state_update_2_port, cyc_state_update_1_port
      , cyc_state_update_0_port, fb_prime_7_port, fb_prime_6_port, 
      fb_prime_5_port, fb_prime_4_port, fb_prime_3_port, fb_prime_2_port, 
      fb_prime_1_port, fb_prime_0_port, plane_2_input_127_port, 
      plane_2_input_126_port, plane_2_input_125_port, plane_2_input_124_port, 
      plane_2_input_123_port, plane_2_input_122_port, plane_2_input_121_port, 
      plane_2_input_120_port, plane_2_input_119_port, plane_2_input_118_port, 
      plane_2_input_117_port, plane_2_input_116_port, plane_2_input_115_port, 
      plane_2_input_114_port, plane_2_input_113_port, plane_2_input_112_port, 
      plane_2_input_111_port, plane_2_input_110_port, plane_2_input_109_port, 
      plane_2_input_108_port, plane_2_input_107_port, plane_2_input_106_port, 
      plane_2_input_105_port, plane_2_input_104_port, plane_2_input_103_port, 
      plane_2_input_102_port, plane_2_input_101_port, plane_2_input_100_port, 
      plane_2_input_99_port, plane_2_input_98_port, plane_2_input_97_port, 
      plane_2_input_96_port, plane_2_input_95_port, plane_2_input_94_port, 
      plane_2_input_93_port, plane_2_input_92_port, plane_2_input_91_port, 
      plane_2_input_90_port, plane_2_input_89_port, plane_2_input_88_port, 
      plane_2_input_87_port, plane_2_input_86_port, plane_2_input_85_port, 
      plane_2_input_84_port, plane_2_input_83_port, plane_2_input_82_port, 
      plane_2_input_81_port, plane_2_input_80_port, plane_2_input_79_port, 
      plane_2_input_78_port, plane_2_input_77_port, plane_2_input_76_port, 
      plane_2_input_75_port, plane_2_input_74_port, plane_2_input_73_port, 
      plane_2_input_72_port, plane_2_input_71_port, plane_2_input_70_port, 
      plane_2_input_69_port, plane_2_input_68_port, plane_2_input_67_port, 
      plane_2_input_66_port, plane_2_input_65_port, plane_2_input_64_port, 
      plane_2_input_63_port, plane_2_input_62_port, plane_2_input_61_port, 
      plane_2_input_60_port, plane_2_input_59_port, plane_2_input_58_port, 
      plane_2_input_57_port, plane_2_input_56_port, plane_2_input_55_port, 
      plane_2_input_54_port, plane_2_input_53_port, plane_2_input_52_port, 
      plane_2_input_51_port, plane_2_input_50_port, plane_2_input_49_port, 
      plane_2_input_48_port, plane_2_input_47_port, plane_2_input_46_port, 
      plane_2_input_45_port, plane_2_input_44_port, plane_2_input_43_port, 
      plane_2_input_42_port, plane_2_input_41_port, plane_2_input_40_port, 
      plane_2_input_39_port, plane_2_input_38_port, plane_2_input_37_port, 
      plane_2_input_36_port, plane_2_input_35_port, plane_2_input_34_port, 
      plane_2_input_33_port, plane_2_input_32_port, plane_2_input_23, 
      plane_2_input_22, plane_2_input_21, plane_2_input_20, plane_2_input_19, 
      plane_2_input_18, plane_2_input_17, plane_2_input_16, plane_2_input_15, 
      plane_2_input_14, plane_2_input_13, plane_2_input_12, plane_2_input_11, 
      plane_2_input_10, plane_2_input_9, plane_2_input_8, plane_2_input_7, 
      plane_2_input_6, plane_2_input_5, plane_2_input_4, plane_2_input_3, 
      plane_2_input_2, plane_2_input_1, plane_2_input_0, N181, N182, 
      state_main_in_p0_127_port, state_main_in_p0_126_port, 
      state_main_in_p0_125_port, state_main_in_p0_124_port, 
      state_main_in_p0_123_port, state_main_in_p0_122_port, 
      state_main_in_p0_121_port, state_main_in_p0_120_port, 
      state_main_in_p0_119_port, state_main_in_p0_118_port, 
      state_main_in_p0_117_port, state_main_in_p0_116_port, 
      state_main_in_p0_115_port, state_main_in_p0_114_port, 
      state_main_in_p0_113_port, state_main_in_p0_112_port, 
      state_main_in_p0_111_port, state_main_in_p0_110_port, 
      state_main_in_p0_109_port, state_main_in_p0_108_port, 
      state_main_in_p0_107_port, state_main_in_p0_106_port, 
      state_main_in_p0_105_port, state_main_in_p0_104_port, 
      state_main_in_p0_103_port, state_main_in_p0_102_port, 
      state_main_in_p0_101_port, state_main_in_p0_100_port, 
      state_main_in_p0_99_port, state_main_in_p0_98_port, 
      state_main_in_p0_97_port, state_main_in_p0_96_port, 
      state_main_in_p0_95_port, state_main_in_p0_94_port, 
      state_main_in_p0_93_port, state_main_in_p0_92_port, 
      state_main_in_p0_91_port, state_main_in_p0_90_port, 
      state_main_in_p0_89_port, state_main_in_p0_88_port, 
      state_main_in_p0_87_port, state_main_in_p0_86_port, 
      state_main_in_p0_85_port, state_main_in_p0_84_port, 
      state_main_in_p0_83_port, state_main_in_p0_82_port, 
      state_main_in_p0_81_port, state_main_in_p0_80_port, 
      state_main_in_p0_79_port, state_main_in_p0_78_port, 
      state_main_in_p0_77_port, state_main_in_p0_76_port, 
      state_main_in_p0_75_port, state_main_in_p0_74_port, 
      state_main_in_p0_73_port, state_main_in_p0_72_port, 
      state_main_in_p0_71_port, state_main_in_p0_70_port, 
      state_main_in_p0_69_port, state_main_in_p0_68_port, 
      state_main_in_p0_67_port, state_main_in_p0_66_port, 
      state_main_in_p0_65_port, state_main_in_p0_64_port, 
      state_main_in_p0_63_port, state_main_in_p0_62_port, 
      state_main_in_p0_61_port, state_main_in_p0_60_port, 
      state_main_in_p0_59_port, state_main_in_p0_58_port, 
      state_main_in_p0_57_port, state_main_in_p0_56_port, 
      state_main_in_p0_55_port, state_main_in_p0_54_port, 
      state_main_in_p0_53_port, state_main_in_p0_52_port, 
      state_main_in_p0_51_port, state_main_in_p0_50_port, 
      state_main_in_p0_49_port, state_main_in_p0_48_port, 
      state_main_in_p0_47_port, state_main_in_p0_46_port, 
      state_main_in_p0_45_port, state_main_in_p0_44_port, 
      state_main_in_p0_43_port, state_main_in_p0_42_port, 
      state_main_in_p0_41_port, state_main_in_p0_40_port, 
      state_main_in_p0_39_port, state_main_in_p0_38_port, 
      state_main_in_p0_37_port, state_main_in_p0_36_port, 
      state_main_in_p0_35_port, state_main_in_p0_34_port, 
      state_main_in_p0_33_port, state_main_in_p0_32_port, 
      state_main_in_p0_31_port, state_main_in_p0_30_port, 
      state_main_in_p0_29_port, state_main_in_p0_28_port, 
      state_main_in_p0_27_port, state_main_in_p0_26_port, 
      state_main_in_p0_25_port, state_main_in_p0_24_port, 
      state_main_in_p0_23_port, state_main_in_p0_22_port, 
      state_main_in_p0_21_port, state_main_in_p0_20_port, 
      state_main_in_p0_19_port, state_main_in_p0_18_port, 
      state_main_in_p0_17_port, state_main_in_p0_16_port, 
      state_main_in_p0_15_port, state_main_in_p0_14_port, 
      state_main_in_p0_13_port, state_main_in_p0_12_port, 
      state_main_in_p0_11_port, state_main_in_p0_10_port, 
      state_main_in_p0_9_port, state_main_in_p0_8_port, state_main_in_p0_7_port
      , state_main_in_p0_6_port, state_main_in_p0_5_port, 
      state_main_in_p0_4_port, state_main_in_p0_3_port, state_main_in_p0_2_port
      , state_main_in_p0_1_port, state_main_in_p0_0_port, perm_output_383_port,
      perm_output_382_port, perm_output_381_port, perm_output_380_port, 
      perm_output_379_port, perm_output_378_port, perm_output_377_port, 
      perm_output_376_port, perm_output_375_port, perm_output_374_port, 
      perm_output_373_port, perm_output_372_port, perm_output_371_port, 
      perm_output_370_port, perm_output_369_port, perm_output_368_port, 
      perm_output_367_port, perm_output_366_port, perm_output_365_port, 
      perm_output_364_port, perm_output_363_port, perm_output_362_port, 
      perm_output_361_port, perm_output_360_port, perm_output_359_port, 
      perm_output_358_port, perm_output_357_port, perm_output_356_port, 
      perm_output_355_port, perm_output_354_port, perm_output_353_port, 
      perm_output_352_port, perm_output_351_port, perm_output_350_port, 
      perm_output_349_port, perm_output_348_port, perm_output_347_port, 
      perm_output_346_port, perm_output_345_port, perm_output_344_port, 
      perm_output_343_port, perm_output_342_port, perm_output_341_port, 
      perm_output_340_port, perm_output_339_port, perm_output_338_port, 
      perm_output_337_port, perm_output_336_port, perm_output_335_port, 
      perm_output_334_port, perm_output_333_port, perm_output_332_port, 
      perm_output_331_port, perm_output_330_port, perm_output_329_port, 
      perm_output_328_port, perm_output_327_port, perm_output_326_port, 
      perm_output_325_port, perm_output_324_port, perm_output_323_port, 
      perm_output_322_port, perm_output_321_port, perm_output_320_port, 
      perm_output_319_port, perm_output_318_port, perm_output_317_port, 
      perm_output_316_port, perm_output_315_port, perm_output_314_port, 
      perm_output_313_port, perm_output_312_port, perm_output_311_port, 
      perm_output_310_port, perm_output_309_port, perm_output_308_port, 
      perm_output_307_port, perm_output_306_port, perm_output_305_port, 
      perm_output_304_port, perm_output_303_port, perm_output_302_port, 
      perm_output_301_port, perm_output_300_port, perm_output_299_port, 
      perm_output_298_port, perm_output_297_port, perm_output_296_port, 
      perm_output_295_port, perm_output_294_port, perm_output_293_port, 
      perm_output_292_port, perm_output_291_port, perm_output_290_port, 
      perm_output_289_port, perm_output_288_port, perm_output_287_port, 
      perm_output_286_port, perm_output_285_port, perm_output_284_port, 
      perm_output_283_port, perm_output_282_port, perm_output_281_port, 
      perm_output_280_port, perm_output_279_port, perm_output_278_port, 
      perm_output_277_port, perm_output_276_port, perm_output_275_port, 
      perm_output_274_port, perm_output_273_port, perm_output_272_port, 
      perm_output_271_port, perm_output_270_port, perm_output_269_port, 
      perm_output_268_port, perm_output_267_port, perm_output_266_port, 
      perm_output_265_port, perm_output_264_port, perm_output_263_port, 
      perm_output_262_port, perm_output_261_port, perm_output_260_port, 
      perm_output_259_port, perm_output_258_port, perm_output_257_port, 
      perm_output_256_port, perm_output_255_port, perm_output_254_port, 
      perm_output_253_port, perm_output_252_port, perm_output_251_port, 
      perm_output_250_port, perm_output_249_port, perm_output_248_port, 
      perm_output_247_port, perm_output_246_port, perm_output_245_port, 
      perm_output_244_port, perm_output_243_port, perm_output_242_port, 
      perm_output_241_port, perm_output_240_port, perm_output_239_port, 
      perm_output_238_port, perm_output_237_port, perm_output_236_port, 
      perm_output_235_port, perm_output_234_port, perm_output_233_port, 
      perm_output_232_port, perm_output_231_port, perm_output_230_port, 
      perm_output_229_port, perm_output_228_port, perm_output_227_port, 
      perm_output_226_port, perm_output_225_port, perm_output_224_port, 
      perm_output_223_port, perm_output_222_port, perm_output_221_port, 
      perm_output_220_port, perm_output_219_port, perm_output_218_port, 
      perm_output_217_port, perm_output_216_port, perm_output_215_port, 
      perm_output_214_port, perm_output_213_port, perm_output_212_port, 
      perm_output_211_port, perm_output_210_port, perm_output_209_port, 
      perm_output_208_port, perm_output_207_port, perm_output_206_port, 
      perm_output_205_port, perm_output_204_port, perm_output_203_port, 
      perm_output_202_port, perm_output_201_port, perm_output_200_port, 
      perm_output_199_port, perm_output_198_port, perm_output_197_port, 
      perm_output_196_port, perm_output_195_port, perm_output_194_port, 
      perm_output_193_port, perm_output_192_port, perm_output_191_port, 
      perm_output_190_port, perm_output_189_port, perm_output_188_port, 
      perm_output_187_port, perm_output_186_port, perm_output_185_port, 
      perm_output_184_port, perm_output_183_port, perm_output_182_port, 
      perm_output_181_port, perm_output_180_port, perm_output_179_port, 
      perm_output_178_port, perm_output_177_port, perm_output_176_port, 
      perm_output_175_port, perm_output_174_port, perm_output_173_port, 
      perm_output_172_port, perm_output_171_port, perm_output_170_port, 
      perm_output_169_port, perm_output_168_port, perm_output_167_port, 
      perm_output_166_port, perm_output_165_port, perm_output_164_port, 
      perm_output_163_port, perm_output_162_port, perm_output_161_port, 
      perm_output_160_port, perm_output_159_port, perm_output_158_port, 
      perm_output_157_port, perm_output_156_port, perm_output_155_port, 
      perm_output_154_port, perm_output_153_port, perm_output_152_port, 
      perm_output_151_port, perm_output_150_port, perm_output_149_port, 
      perm_output_148_port, perm_output_147_port, perm_output_146_port, 
      perm_output_145_port, perm_output_144_port, perm_output_143_port, 
      perm_output_142_port, perm_output_141_port, perm_output_140_port, 
      perm_output_139_port, perm_output_138_port, perm_output_137_port, 
      perm_output_136_port, perm_output_135_port, perm_output_134_port, 
      perm_output_133_port, perm_output_132_port, perm_output_131_port, 
      perm_output_130_port, perm_output_129_port, perm_output_128_port, 
      perm_output_127_port, perm_output_126_port, perm_output_125_port, 
      perm_output_124_port, perm_output_123_port, perm_output_122_port, 
      perm_output_121_port, perm_output_120_port, perm_output_119_port, 
      perm_output_118_port, perm_output_117_port, perm_output_116_port, 
      perm_output_115_port, perm_output_114_port, perm_output_113_port, 
      perm_output_112_port, perm_output_111_port, perm_output_110_port, 
      perm_output_109_port, perm_output_108_port, perm_output_107_port, 
      perm_output_106_port, perm_output_105_port, perm_output_104_port, 
      perm_output_103_port, perm_output_102_port, perm_output_101_port, 
      perm_output_100_port, perm_output_99_port, perm_output_98_port, 
      perm_output_97_port, perm_output_96_port, perm_output_95_port, 
      perm_output_94_port, perm_output_93_port, perm_output_92_port, 
      perm_output_91_port, perm_output_90_port, perm_output_89_port, 
      perm_output_88_port, perm_output_87_port, perm_output_86_port, 
      perm_output_85_port, perm_output_84_port, perm_output_83_port, 
      perm_output_82_port, perm_output_81_port, perm_output_80_port, 
      perm_output_79_port, perm_output_78_port, perm_output_77_port, 
      perm_output_76_port, perm_output_75_port, perm_output_74_port, 
      perm_output_73_port, perm_output_72_port, perm_output_71_port, 
      perm_output_70_port, perm_output_69_port, perm_output_68_port, 
      perm_output_67_port, perm_output_66_port, perm_output_65_port, 
      perm_output_64_port, perm_output_63_port, perm_output_62_port, 
      perm_output_61_port, perm_output_60_port, perm_output_59_port, 
      perm_output_58_port, perm_output_57_port, perm_output_56_port, 
      perm_output_55_port, perm_output_54_port, perm_output_53_port, 
      perm_output_52_port, perm_output_51_port, perm_output_50_port, 
      perm_output_49_port, perm_output_48_port, perm_output_47_port, 
      perm_output_46_port, perm_output_45_port, perm_output_44_port, 
      perm_output_43_port, perm_output_42_port, perm_output_41_port, 
      perm_output_40_port, perm_output_39_port, perm_output_38_port, 
      perm_output_37_port, perm_output_36_port, perm_output_35_port, 
      perm_output_34_port, perm_output_33_port, perm_output_32_port, 
      perm_output_31_port, perm_output_30_port, perm_output_29_port, 
      perm_output_28_port, perm_output_27_port, perm_output_26_port, 
      perm_output_25_port, perm_output_24_port, perm_output_23_port, 
      perm_output_22_port, perm_output_21_port, perm_output_20_port, 
      perm_output_19_port, perm_output_18_port, perm_output_17_port, 
      perm_output_16_port, perm_output_15_port, perm_output_14_port, 
      perm_output_13_port, perm_output_12_port, perm_output_11_port, 
      perm_output_10_port, perm_output_9_port, perm_output_8_port, 
      perm_output_7_port, perm_output_6_port, perm_output_5_port, 
      perm_output_4_port, perm_output_3_port, perm_output_2_port, 
      perm_output_1_port, perm_output_0_port, N183, N184, N185, N186, N187, 
      N188, N189, N190, N191, N192, N193, N194, N195, N196, N197, N198, N199, 
      N200, N201, N202, N203, N204, N205, N206, N207, N208, N209, N210, N211, 
      N212, N213, N214, N215, N216, N217, N218, N219, N220, N221, N222, N223, 
      N224, N225, N226, N227, N228, N229, N230, N231, N232, N233, N234, N235, 
      N236, N237, N238, N239, N240, N241, N242, N243, N244, N245, N246, N247, 
      N248, N249, N250, N251, N252, N253, N254, N255, N256, N257, N258, N259, 
      N260, N261, N262, N263, N264, N265, N266, N267, N268, N269, N270, N271, 
      N272, N273, N274, N275, N276, N277, N278, N279, N280, N281, N282, N283, 
      N284, N285, N286, N287, N288, N289, N290, N291, N292, N293, N294, N295, 
      N296, N297, N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, 
      N308, N309, N310, N311, N312, state_main_in_p1_127_port, 
      state_main_in_p1_126_port, state_main_in_p1_125_port, 
      state_main_in_p1_124_port, state_main_in_p1_123_port, 
      state_main_in_p1_122_port, state_main_in_p1_121_port, 
      state_main_in_p1_120_port, state_main_in_p1_119_port, 
      state_main_in_p1_118_port, state_main_in_p1_117_port, 
      state_main_in_p1_116_port, state_main_in_p1_115_port, 
      state_main_in_p1_114_port, state_main_in_p1_113_port, 
      state_main_in_p1_112_port, state_main_in_p1_111_port, 
      state_main_in_p1_110_port, state_main_in_p1_109_port, 
      state_main_in_p1_108_port, state_main_in_p1_107_port, 
      state_main_in_p1_106_port, state_main_in_p1_105_port, 
      state_main_in_p1_104_port, state_main_in_p1_103_port, 
      state_main_in_p1_102_port, state_main_in_p1_101_port, 
      state_main_in_p1_100_port, state_main_in_p1_99_port, 
      state_main_in_p1_98_port, state_main_in_p1_97_port, 
      state_main_in_p1_96_port, state_main_in_p1_95_port, 
      state_main_in_p1_94_port, state_main_in_p1_93_port, 
      state_main_in_p1_92_port, state_main_in_p1_91_port, 
      state_main_in_p1_90_port, state_main_in_p1_89_port, 
      state_main_in_p1_88_port, state_main_in_p1_87_port, 
      state_main_in_p1_86_port, state_main_in_p1_85_port, 
      state_main_in_p1_84_port, state_main_in_p1_83_port, 
      state_main_in_p1_82_port, state_main_in_p1_81_port, 
      state_main_in_p1_80_port, state_main_in_p1_79_port, 
      state_main_in_p1_78_port, state_main_in_p1_77_port, 
      state_main_in_p1_76_port, state_main_in_p1_75_port, 
      state_main_in_p1_74_port, state_main_in_p1_73_port, 
      state_main_in_p1_72_port, state_main_in_p1_71_port, 
      state_main_in_p1_70_port, state_main_in_p1_69_port, 
      state_main_in_p1_68_port, state_main_in_p1_67_port, 
      state_main_in_p1_66_port, state_main_in_p1_65_port, 
      state_main_in_p1_64_port, state_main_in_p1_63_port, 
      state_main_in_p1_62_port, state_main_in_p1_61_port, 
      state_main_in_p1_60_port, state_main_in_p1_59_port, 
      state_main_in_p1_58_port, state_main_in_p1_57_port, 
      state_main_in_p1_56_port, state_main_in_p1_55_port, 
      state_main_in_p1_54_port, state_main_in_p1_53_port, 
      state_main_in_p1_52_port, state_main_in_p1_51_port, 
      state_main_in_p1_50_port, state_main_in_p1_49_port, 
      state_main_in_p1_48_port, state_main_in_p1_47_port, 
      state_main_in_p1_46_port, state_main_in_p1_45_port, 
      state_main_in_p1_44_port, state_main_in_p1_43_port, 
      state_main_in_p1_42_port, state_main_in_p1_41_port, 
      state_main_in_p1_40_port, state_main_in_p1_39_port, 
      state_main_in_p1_38_port, state_main_in_p1_37_port, 
      state_main_in_p1_36_port, state_main_in_p1_35_port, 
      state_main_in_p1_34_port, state_main_in_p1_33_port, 
      state_main_in_p1_32_port, state_main_in_p1_31_port, 
      state_main_in_p1_30_port, state_main_in_p1_29_port, 
      state_main_in_p1_28_port, state_main_in_p1_27_port, 
      state_main_in_p1_26_port, state_main_in_p1_25_port, 
      state_main_in_p1_24_port, state_main_in_p1_23_port, 
      state_main_in_p1_22_port, state_main_in_p1_21_port, 
      state_main_in_p1_20_port, state_main_in_p1_19_port, 
      state_main_in_p1_18_port, state_main_in_p1_17_port, 
      state_main_in_p1_16_port, state_main_in_p1_15_port, 
      state_main_in_p1_14_port, state_main_in_p1_13_port, 
      state_main_in_p1_12_port, state_main_in_p1_11_port, 
      state_main_in_p1_10_port, state_main_in_p1_9_port, 
      state_main_in_p1_8_port, state_main_in_p1_7_port, state_main_in_p1_6_port
      , state_main_in_p1_5_port, state_main_in_p1_4_port, 
      state_main_in_p1_3_port, state_main_in_p1_2_port, state_main_in_p1_1_port
      , state_main_in_p1_0_port, N313, N314, N315, N316, N317, N318, N319, N320
      , N321, N322, N323, N324, N325, N326, N327, N328, N329, N330, N331, N332,
      N333, N334, N335, N336, N337, N338, N339, N340, N341, N342, N343, N344, 
      N345, N346, N347, N348, N349, N350, N351, N352, N353, N354, N355, N356, 
      N357, N358, N359, N360, N361, N362, N363, N364, N365, N366, N367, N368, 
      N369, N370, N371, N372, N373, N374, N375, N376, N377, N378, N379, N380, 
      N381, N382, N383, N384, N385, N386, N387, N388, N389, N390, N391, N392, 
      N393, N394, N395, N396, N397, N398, N399, N400, N401, N402, N403, N404, 
      N405, N406, N407, N408, N409, N410, N411, N412, N413, N414, N415, N416, 
      N417, N418, N419, N420, N421, N422, N423, N424, N425, N426, N427, N428, 
      N429, N430, N431, N432, N433, N434, N435, N436, N437, N438, N439, N440, 
      N441, N442, state_main_in_p2_127_port, state_main_in_p2_126_port, 
      state_main_in_p2_125_port, state_main_in_p2_124_port, 
      state_main_in_p2_123_port, state_main_in_p2_122_port, 
      state_main_in_p2_121_port, state_main_in_p2_120_port, 
      state_main_in_p2_119_port, state_main_in_p2_118_port, 
      state_main_in_p2_117_port, state_main_in_p2_116_port, 
      state_main_in_p2_115_port, state_main_in_p2_114_port, 
      state_main_in_p2_113_port, state_main_in_p2_112_port, 
      state_main_in_p2_111_port, state_main_in_p2_110_port, 
      state_main_in_p2_109_port, state_main_in_p2_108_port, 
      state_main_in_p2_107_port, state_main_in_p2_106_port, 
      state_main_in_p2_105_port, state_main_in_p2_104_port, 
      state_main_in_p2_103_port, state_main_in_p2_102_port, 
      state_main_in_p2_101_port, state_main_in_p2_100_port, 
      state_main_in_p2_99_port, state_main_in_p2_98_port, 
      state_main_in_p2_97_port, state_main_in_p2_96_port, 
      state_main_in_p2_95_port, state_main_in_p2_94_port, 
      state_main_in_p2_93_port, state_main_in_p2_92_port, 
      state_main_in_p2_91_port, state_main_in_p2_90_port, 
      state_main_in_p2_89_port, state_main_in_p2_88_port, 
      state_main_in_p2_87_port, state_main_in_p2_86_port, 
      state_main_in_p2_85_port, state_main_in_p2_84_port, 
      state_main_in_p2_83_port, state_main_in_p2_82_port, 
      state_main_in_p2_81_port, state_main_in_p2_80_port, 
      state_main_in_p2_79_port, state_main_in_p2_78_port, 
      state_main_in_p2_77_port, state_main_in_p2_76_port, 
      state_main_in_p2_75_port, state_main_in_p2_74_port, 
      state_main_in_p2_73_port, state_main_in_p2_72_port, 
      state_main_in_p2_71_port, state_main_in_p2_70_port, 
      state_main_in_p2_69_port, state_main_in_p2_68_port, 
      state_main_in_p2_67_port, state_main_in_p2_66_port, 
      state_main_in_p2_65_port, state_main_in_p2_64_port, 
      state_main_in_p2_63_port, state_main_in_p2_62_port, 
      state_main_in_p2_61_port, state_main_in_p2_60_port, 
      state_main_in_p2_59_port, state_main_in_p2_58_port, 
      state_main_in_p2_57_port, state_main_in_p2_56_port, 
      state_main_in_p2_55_port, state_main_in_p2_54_port, 
      state_main_in_p2_53_port, state_main_in_p2_52_port, 
      state_main_in_p2_51_port, state_main_in_p2_50_port, 
      state_main_in_p2_49_port, state_main_in_p2_48_port, 
      state_main_in_p2_47_port, state_main_in_p2_46_port, 
      state_main_in_p2_45_port, state_main_in_p2_44_port, 
      state_main_in_p2_43_port, state_main_in_p2_42_port, 
      state_main_in_p2_41_port, state_main_in_p2_40_port, 
      state_main_in_p2_39_port, state_main_in_p2_38_port, 
      state_main_in_p2_37_port, state_main_in_p2_36_port, 
      state_main_in_p2_35_port, state_main_in_p2_34_port, 
      state_main_in_p2_33_port, state_main_in_p2_32_port, 
      state_main_in_p2_31_port, state_main_in_p2_30_port, 
      state_main_in_p2_29_port, state_main_in_p2_28_port, 
      state_main_in_p2_27_port, state_main_in_p2_26_port, 
      state_main_in_p2_25_port, state_main_in_p2_24_port, 
      state_main_in_p2_23_port, state_main_in_p2_22_port, 
      state_main_in_p2_21_port, state_main_in_p2_20_port, 
      state_main_in_p2_19_port, state_main_in_p2_18_port, 
      state_main_in_p2_17_port, state_main_in_p2_16_port, 
      state_main_in_p2_15_port, state_main_in_p2_14_port, 
      state_main_in_p2_13_port, state_main_in_p2_12_port, 
      state_main_in_p2_11_port, state_main_in_p2_10_port, 
      state_main_in_p2_9_port, state_main_in_p2_8_port, state_main_in_p2_7_port
      , state_main_in_p2_6_port, state_main_in_p2_5_port, 
      state_main_in_p2_4_port, state_main_in_p2_3_port, state_main_in_p2_2_port
      , state_main_in_p2_1_port, state_main_in_p2_0_port, N443, N444, N445, 
      N446, N447, N448, N449, N450, N451, N452, N453, N454, N455, N456, N457, 
      N458, N459, N460, N461, N462, N463, N464, N465, N466, N467, N468, N469, 
      N470, N471, N472, N473, N474, N475, N476, N477, N478, N479, N480, N481, 
      N482, N483, N484, N485, N486, N487, N488, N489, N490, N491, N492, N493, 
      N494, N495, N496, N497, N498, N499, N500, N501, N502, N503, N504, N505, 
      N506, N507, N508, N509, N510, N511, N512, N513, N514, N515, N516, N517, 
      N518, N519, N520, N521, N522, N523, N524, N525, N526, N527, N528, N529, 
      N530, N531, N532, N533, N534, N535, N536, N537, N538, N539, N540, N541, 
      N542, N543, N544, N545, N546, N547, N548, N549, N550, N551, N552, N553, 
      N554, N555, N556, N557, N558, N559, N560, N561, N562, N563, N564, N565, 
      N566, N567, N568, N569, N570, N571, N572, N573, N574 : std_logic;

begin
   ( bdi_key_31_port, bdi_key_30_port, bdi_key_29_port, bdi_key_28_port, 
      bdi_key_27_port, bdi_key_26_port, bdi_key_25_port, bdi_key_24_port, 
      bdi_key_23_port, bdi_key_22_port, bdi_key_21_port, bdi_key_20_port, 
      bdi_key_19_port, bdi_key_18_port, bdi_key_17_port, bdi_key_16_port, 
      bdi_key_15_port, bdi_key_14_port, bdi_key_13_port, bdi_key_12_port, 
      bdi_key_11_port, bdi_key_10_port, bdi_key_9_port, bdi_key_8_port, 
      bdi_key_7_port, bdi_key_6_port, bdi_key_5_port, bdi_key_4_port, 
      bdi_key_3_port, bdi_key_2_port, bdi_key_1_port, bdi_key_0_port ) <= 
      bdi_key;
   bdo_out <= ( bdo_out_31_port, bdo_out_30_port, bdo_out_29_port, 
      bdo_out_28_port, bdo_out_27_port, bdo_out_26_port, bdo_out_25_port, 
      bdo_out_24_port, bdo_out_23_port, bdo_out_22_port, bdo_out_21_port, 
      bdo_out_20_port, bdo_out_19_port, bdo_out_18_port, bdo_out_17_port, 
      bdo_out_16_port, bdo_out_15_port, bdo_out_14_port, bdo_out_13_port, 
      bdo_out_12_port, bdo_out_11_port, bdo_out_10_port, bdo_out_9_port, 
      bdo_out_8_port, bdo_out_7_port, bdo_out_6_port, bdo_out_5_port, 
      bdo_out_4_port, bdo_out_3_port, bdo_out_2_port, bdo_out_1_port, 
      bdo_out_0_port );
   
   C271 : GTECH_OR2 port map( A => cycd_sel(1), B => N168, Z => N162);
   C274 : GTECH_OR2 port map( A => N167, B => cycd_sel(0), Z => N164);
   C276 : GTECH_AND2 port map( A => cycd_sel(1), B => cycd_sel(0), Z => N166);
   C279 : GTECH_AND2 port map( A => N167, B => N168, Z => N169);
   C421 : GTECH_AND2 port map( A => N170, B => N171, Z => N172);
   C423 : GTECH_OR2 port map( A => dcount_in(1), B => N171, Z => N173);
   C426 : GTECH_OR2 port map( A => N170, B => dcount_in(0), Z => N175);
   C428 : GTECH_AND2 port map( A => dcount_in(1), B => dcount_in(0), Z => N177)
                           ;
   state_main_p0 : reg_custom_LEN128_1 port map( clk => clk, en => 
                           state_main_en(0), din(127) => 
                           state_main_in_p0_127_port, din(126) => 
                           state_main_in_p0_126_port, din(125) => 
                           state_main_in_p0_125_port, din(124) => 
                           state_main_in_p0_124_port, din(123) => 
                           state_main_in_p0_123_port, din(122) => 
                           state_main_in_p0_122_port, din(121) => 
                           state_main_in_p0_121_port, din(120) => 
                           state_main_in_p0_120_port, din(119) => 
                           state_main_in_p0_119_port, din(118) => 
                           state_main_in_p0_118_port, din(117) => 
                           state_main_in_p0_117_port, din(116) => 
                           state_main_in_p0_116_port, din(115) => 
                           state_main_in_p0_115_port, din(114) => 
                           state_main_in_p0_114_port, din(113) => 
                           state_main_in_p0_113_port, din(112) => 
                           state_main_in_p0_112_port, din(111) => 
                           state_main_in_p0_111_port, din(110) => 
                           state_main_in_p0_110_port, din(109) => 
                           state_main_in_p0_109_port, din(108) => 
                           state_main_in_p0_108_port, din(107) => 
                           state_main_in_p0_107_port, din(106) => 
                           state_main_in_p0_106_port, din(105) => 
                           state_main_in_p0_105_port, din(104) => 
                           state_main_in_p0_104_port, din(103) => 
                           state_main_in_p0_103_port, din(102) => 
                           state_main_in_p0_102_port, din(101) => 
                           state_main_in_p0_101_port, din(100) => 
                           state_main_in_p0_100_port, din(99) => 
                           state_main_in_p0_99_port, din(98) => 
                           state_main_in_p0_98_port, din(97) => 
                           state_main_in_p0_97_port, din(96) => 
                           state_main_in_p0_96_port, din(95) => 
                           state_main_in_p0_95_port, din(94) => 
                           state_main_in_p0_94_port, din(93) => 
                           state_main_in_p0_93_port, din(92) => 
                           state_main_in_p0_92_port, din(91) => 
                           state_main_in_p0_91_port, din(90) => 
                           state_main_in_p0_90_port, din(89) => 
                           state_main_in_p0_89_port, din(88) => 
                           state_main_in_p0_88_port, din(87) => 
                           state_main_in_p0_87_port, din(86) => 
                           state_main_in_p0_86_port, din(85) => 
                           state_main_in_p0_85_port, din(84) => 
                           state_main_in_p0_84_port, din(83) => 
                           state_main_in_p0_83_port, din(82) => 
                           state_main_in_p0_82_port, din(81) => 
                           state_main_in_p0_81_port, din(80) => 
                           state_main_in_p0_80_port, din(79) => 
                           state_main_in_p0_79_port, din(78) => 
                           state_main_in_p0_78_port, din(77) => 
                           state_main_in_p0_77_port, din(76) => 
                           state_main_in_p0_76_port, din(75) => 
                           state_main_in_p0_75_port, din(74) => 
                           state_main_in_p0_74_port, din(73) => 
                           state_main_in_p0_73_port, din(72) => 
                           state_main_in_p0_72_port, din(71) => 
                           state_main_in_p0_71_port, din(70) => 
                           state_main_in_p0_70_port, din(69) => 
                           state_main_in_p0_69_port, din(68) => 
                           state_main_in_p0_68_port, din(67) => 
                           state_main_in_p0_67_port, din(66) => 
                           state_main_in_p0_66_port, din(65) => 
                           state_main_in_p0_65_port, din(64) => 
                           state_main_in_p0_64_port, din(63) => 
                           state_main_in_p0_63_port, din(62) => 
                           state_main_in_p0_62_port, din(61) => 
                           state_main_in_p0_61_port, din(60) => 
                           state_main_in_p0_60_port, din(59) => 
                           state_main_in_p0_59_port, din(58) => 
                           state_main_in_p0_58_port, din(57) => 
                           state_main_in_p0_57_port, din(56) => 
                           state_main_in_p0_56_port, din(55) => 
                           state_main_in_p0_55_port, din(54) => 
                           state_main_in_p0_54_port, din(53) => 
                           state_main_in_p0_53_port, din(52) => 
                           state_main_in_p0_52_port, din(51) => 
                           state_main_in_p0_51_port, din(50) => 
                           state_main_in_p0_50_port, din(49) => 
                           state_main_in_p0_49_port, din(48) => 
                           state_main_in_p0_48_port, din(47) => 
                           state_main_in_p0_47_port, din(46) => 
                           state_main_in_p0_46_port, din(45) => 
                           state_main_in_p0_45_port, din(44) => 
                           state_main_in_p0_44_port, din(43) => 
                           state_main_in_p0_43_port, din(42) => 
                           state_main_in_p0_42_port, din(41) => 
                           state_main_in_p0_41_port, din(40) => 
                           state_main_in_p0_40_port, din(39) => 
                           state_main_in_p0_39_port, din(38) => 
                           state_main_in_p0_38_port, din(37) => 
                           state_main_in_p0_37_port, din(36) => 
                           state_main_in_p0_36_port, din(35) => 
                           state_main_in_p0_35_port, din(34) => 
                           state_main_in_p0_34_port, din(33) => 
                           state_main_in_p0_33_port, din(32) => 
                           state_main_in_p0_32_port, din(31) => 
                           state_main_in_p0_31_port, din(30) => 
                           state_main_in_p0_30_port, din(29) => 
                           state_main_in_p0_29_port, din(28) => 
                           state_main_in_p0_28_port, din(27) => 
                           state_main_in_p0_27_port, din(26) => 
                           state_main_in_p0_26_port, din(25) => 
                           state_main_in_p0_25_port, din(24) => 
                           state_main_in_p0_24_port, din(23) => 
                           state_main_in_p0_23_port, din(22) => 
                           state_main_in_p0_22_port, din(21) => 
                           state_main_in_p0_21_port, din(20) => 
                           state_main_in_p0_20_port, din(19) => 
                           state_main_in_p0_19_port, din(18) => 
                           state_main_in_p0_18_port, din(17) => 
                           state_main_in_p0_17_port, din(16) => 
                           state_main_in_p0_16_port, din(15) => 
                           state_main_in_p0_15_port, din(14) => 
                           state_main_in_p0_14_port, din(13) => 
                           state_main_in_p0_13_port, din(12) => 
                           state_main_in_p0_12_port, din(11) => 
                           state_main_in_p0_11_port, din(10) => 
                           state_main_in_p0_10_port, din(9) => 
                           state_main_in_p0_9_port, din(8) => 
                           state_main_in_p0_8_port, din(7) => 
                           state_main_in_p0_7_port, din(6) => 
                           state_main_in_p0_6_port, din(5) => 
                           state_main_in_p0_5_port, din(4) => 
                           state_main_in_p0_4_port, din(3) => 
                           state_main_in_p0_3_port, din(2) => 
                           state_main_in_p0_2_port, din(1) => 
                           state_main_in_p0_1_port, din(0) => 
                           state_main_in_p0_0_port, qout(127) => 
                           state_main_out_plane0_127_port, qout(126) => 
                           state_main_out_plane0_126_port, qout(125) => 
                           state_main_out_plane0_125_port, qout(124) => 
                           state_main_out_plane0_124_port, qout(123) => 
                           state_main_out_plane0_123_port, qout(122) => 
                           state_main_out_plane0_122_port, qout(121) => 
                           state_main_out_plane0_121_port, qout(120) => 
                           state_main_out_plane0_120_port, qout(119) => 
                           state_main_out_plane0_119_port, qout(118) => 
                           state_main_out_plane0_118_port, qout(117) => 
                           state_main_out_plane0_117_port, qout(116) => 
                           state_main_out_plane0_116_port, qout(115) => 
                           state_main_out_plane0_115_port, qout(114) => 
                           state_main_out_plane0_114_port, qout(113) => 
                           state_main_out_plane0_113_port, qout(112) => 
                           state_main_out_plane0_112_port, qout(111) => 
                           state_main_out_plane0_111_port, qout(110) => 
                           state_main_out_plane0_110_port, qout(109) => 
                           state_main_out_plane0_109_port, qout(108) => 
                           state_main_out_plane0_108_port, qout(107) => 
                           state_main_out_plane0_107_port, qout(106) => 
                           state_main_out_plane0_106_port, qout(105) => 
                           state_main_out_plane0_105_port, qout(104) => 
                           state_main_out_plane0_104_port, qout(103) => 
                           state_main_out_plane0_103_port, qout(102) => 
                           state_main_out_plane0_102_port, qout(101) => 
                           state_main_out_plane0_101_port, qout(100) => 
                           state_main_out_plane0_100_port, qout(99) => 
                           state_main_out_plane0_99_port, qout(98) => 
                           state_main_out_plane0_98_port, qout(97) => 
                           state_main_out_plane0_97_port, qout(96) => 
                           state_main_out_plane0_96_port, qout(95) => 
                           state_main_out_plane0_95_port, qout(94) => 
                           state_main_out_plane0_94_port, qout(93) => 
                           state_main_out_plane0_93_port, qout(92) => 
                           state_main_out_plane0_92_port, qout(91) => 
                           state_main_out_plane0_91_port, qout(90) => 
                           state_main_out_plane0_90_port, qout(89) => 
                           state_main_out_plane0_89_port, qout(88) => 
                           state_main_out_plane0_88_port, qout(87) => 
                           state_main_out_plane0_87_port, qout(86) => 
                           state_main_out_plane0_86_port, qout(85) => 
                           state_main_out_plane0_85_port, qout(84) => 
                           state_main_out_plane0_84_port, qout(83) => 
                           state_main_out_plane0_83_port, qout(82) => 
                           state_main_out_plane0_82_port, qout(81) => 
                           state_main_out_plane0_81_port, qout(80) => 
                           state_main_out_plane0_80_port, qout(79) => 
                           state_main_out_plane0_79_port, qout(78) => 
                           state_main_out_plane0_78_port, qout(77) => 
                           state_main_out_plane0_77_port, qout(76) => 
                           state_main_out_plane0_76_port, qout(75) => 
                           state_main_out_plane0_75_port, qout(74) => 
                           state_main_out_plane0_74_port, qout(73) => 
                           state_main_out_plane0_73_port, qout(72) => 
                           state_main_out_plane0_72_port, qout(71) => 
                           state_main_out_plane0_71_port, qout(70) => 
                           state_main_out_plane0_70_port, qout(69) => 
                           state_main_out_plane0_69_port, qout(68) => 
                           state_main_out_plane0_68_port, qout(67) => 
                           state_main_out_plane0_67_port, qout(66) => 
                           state_main_out_plane0_66_port, qout(65) => 
                           state_main_out_plane0_65_port, qout(64) => 
                           state_main_out_plane0_64_port, qout(63) => 
                           state_main_out_plane0_63_port, qout(62) => 
                           state_main_out_plane0_62_port, qout(61) => 
                           state_main_out_plane0_61_port, qout(60) => 
                           state_main_out_plane0_60_port, qout(59) => 
                           state_main_out_plane0_59_port, qout(58) => 
                           state_main_out_plane0_58_port, qout(57) => 
                           state_main_out_plane0_57_port, qout(56) => 
                           state_main_out_plane0_56_port, qout(55) => 
                           state_main_out_plane0_55_port, qout(54) => 
                           state_main_out_plane0_54_port, qout(53) => 
                           state_main_out_plane0_53_port, qout(52) => 
                           state_main_out_plane0_52_port, qout(51) => 
                           state_main_out_plane0_51_port, qout(50) => 
                           state_main_out_plane0_50_port, qout(49) => 
                           state_main_out_plane0_49_port, qout(48) => 
                           state_main_out_plane0_48_port, qout(47) => 
                           state_main_out_plane0_47_port, qout(46) => 
                           state_main_out_plane0_46_port, qout(45) => 
                           state_main_out_plane0_45_port, qout(44) => 
                           state_main_out_plane0_44_port, qout(43) => 
                           state_main_out_plane0_43_port, qout(42) => 
                           state_main_out_plane0_42_port, qout(41) => 
                           state_main_out_plane0_41_port, qout(40) => 
                           state_main_out_plane0_40_port, qout(39) => 
                           state_main_out_plane0_39_port, qout(38) => 
                           state_main_out_plane0_38_port, qout(37) => 
                           state_main_out_plane0_37_port, qout(36) => 
                           state_main_out_plane0_36_port, qout(35) => 
                           state_main_out_plane0_35_port, qout(34) => 
                           state_main_out_plane0_34_port, qout(33) => 
                           state_main_out_plane0_33_port, qout(32) => 
                           state_main_out_plane0_32_port, qout(31) => 
                           state_main_out_plane0_31_port, qout(30) => 
                           state_main_out_plane0_30_port, qout(29) => 
                           state_main_out_plane0_29_port, qout(28) => 
                           state_main_out_plane0_28_port, qout(27) => 
                           state_main_out_plane0_27_port, qout(26) => 
                           state_main_out_plane0_26_port, qout(25) => 
                           state_main_out_plane0_25_port, qout(24) => 
                           state_main_out_plane0_24_port, qout(23) => 
                           state_main_out_plane0_23_port, qout(22) => 
                           state_main_out_plane0_22_port, qout(21) => 
                           state_main_out_plane0_21_port, qout(20) => 
                           state_main_out_plane0_20_port, qout(19) => 
                           state_main_out_plane0_19_port, qout(18) => 
                           state_main_out_plane0_18_port, qout(17) => 
                           state_main_out_plane0_17_port, qout(16) => 
                           state_main_out_plane0_16_port, qout(15) => 
                           state_main_out_plane0_15_port, qout(14) => 
                           state_main_out_plane0_14_port, qout(13) => 
                           state_main_out_plane0_13_port, qout(12) => 
                           state_main_out_plane0_12_port, qout(11) => 
                           state_main_out_plane0_11_port, qout(10) => 
                           state_main_out_plane0_10_port, qout(9) => 
                           state_main_out_plane0_9_port, qout(8) => 
                           state_main_out_plane0_8_port, qout(7) => 
                           state_main_out_plane0_7_port, qout(6) => 
                           state_main_out_plane0_6_port, qout(5) => 
                           state_main_out_plane0_5_port, qout(4) => 
                           state_main_out_plane0_4_port, qout(3) => 
                           state_main_out_plane0_3_port, qout(2) => 
                           state_main_out_plane0_2_port, qout(1) => 
                           state_main_out_plane0_1_port, qout(0) => 
                           state_main_out_plane0_0_port);
   state_main_p1 : reg_custom_LEN128_1 port map( clk => clk, en => 
                           state_main_en(1), din(127) => 
                           state_main_in_p1_127_port, din(126) => 
                           state_main_in_p1_126_port, din(125) => 
                           state_main_in_p1_125_port, din(124) => 
                           state_main_in_p1_124_port, din(123) => 
                           state_main_in_p1_123_port, din(122) => 
                           state_main_in_p1_122_port, din(121) => 
                           state_main_in_p1_121_port, din(120) => 
                           state_main_in_p1_120_port, din(119) => 
                           state_main_in_p1_119_port, din(118) => 
                           state_main_in_p1_118_port, din(117) => 
                           state_main_in_p1_117_port, din(116) => 
                           state_main_in_p1_116_port, din(115) => 
                           state_main_in_p1_115_port, din(114) => 
                           state_main_in_p1_114_port, din(113) => 
                           state_main_in_p1_113_port, din(112) => 
                           state_main_in_p1_112_port, din(111) => 
                           state_main_in_p1_111_port, din(110) => 
                           state_main_in_p1_110_port, din(109) => 
                           state_main_in_p1_109_port, din(108) => 
                           state_main_in_p1_108_port, din(107) => 
                           state_main_in_p1_107_port, din(106) => 
                           state_main_in_p1_106_port, din(105) => 
                           state_main_in_p1_105_port, din(104) => 
                           state_main_in_p1_104_port, din(103) => 
                           state_main_in_p1_103_port, din(102) => 
                           state_main_in_p1_102_port, din(101) => 
                           state_main_in_p1_101_port, din(100) => 
                           state_main_in_p1_100_port, din(99) => 
                           state_main_in_p1_99_port, din(98) => 
                           state_main_in_p1_98_port, din(97) => 
                           state_main_in_p1_97_port, din(96) => 
                           state_main_in_p1_96_port, din(95) => 
                           state_main_in_p1_95_port, din(94) => 
                           state_main_in_p1_94_port, din(93) => 
                           state_main_in_p1_93_port, din(92) => 
                           state_main_in_p1_92_port, din(91) => 
                           state_main_in_p1_91_port, din(90) => 
                           state_main_in_p1_90_port, din(89) => 
                           state_main_in_p1_89_port, din(88) => 
                           state_main_in_p1_88_port, din(87) => 
                           state_main_in_p1_87_port, din(86) => 
                           state_main_in_p1_86_port, din(85) => 
                           state_main_in_p1_85_port, din(84) => 
                           state_main_in_p1_84_port, din(83) => 
                           state_main_in_p1_83_port, din(82) => 
                           state_main_in_p1_82_port, din(81) => 
                           state_main_in_p1_81_port, din(80) => 
                           state_main_in_p1_80_port, din(79) => 
                           state_main_in_p1_79_port, din(78) => 
                           state_main_in_p1_78_port, din(77) => 
                           state_main_in_p1_77_port, din(76) => 
                           state_main_in_p1_76_port, din(75) => 
                           state_main_in_p1_75_port, din(74) => 
                           state_main_in_p1_74_port, din(73) => 
                           state_main_in_p1_73_port, din(72) => 
                           state_main_in_p1_72_port, din(71) => 
                           state_main_in_p1_71_port, din(70) => 
                           state_main_in_p1_70_port, din(69) => 
                           state_main_in_p1_69_port, din(68) => 
                           state_main_in_p1_68_port, din(67) => 
                           state_main_in_p1_67_port, din(66) => 
                           state_main_in_p1_66_port, din(65) => 
                           state_main_in_p1_65_port, din(64) => 
                           state_main_in_p1_64_port, din(63) => 
                           state_main_in_p1_63_port, din(62) => 
                           state_main_in_p1_62_port, din(61) => 
                           state_main_in_p1_61_port, din(60) => 
                           state_main_in_p1_60_port, din(59) => 
                           state_main_in_p1_59_port, din(58) => 
                           state_main_in_p1_58_port, din(57) => 
                           state_main_in_p1_57_port, din(56) => 
                           state_main_in_p1_56_port, din(55) => 
                           state_main_in_p1_55_port, din(54) => 
                           state_main_in_p1_54_port, din(53) => 
                           state_main_in_p1_53_port, din(52) => 
                           state_main_in_p1_52_port, din(51) => 
                           state_main_in_p1_51_port, din(50) => 
                           state_main_in_p1_50_port, din(49) => 
                           state_main_in_p1_49_port, din(48) => 
                           state_main_in_p1_48_port, din(47) => 
                           state_main_in_p1_47_port, din(46) => 
                           state_main_in_p1_46_port, din(45) => 
                           state_main_in_p1_45_port, din(44) => 
                           state_main_in_p1_44_port, din(43) => 
                           state_main_in_p1_43_port, din(42) => 
                           state_main_in_p1_42_port, din(41) => 
                           state_main_in_p1_41_port, din(40) => 
                           state_main_in_p1_40_port, din(39) => 
                           state_main_in_p1_39_port, din(38) => 
                           state_main_in_p1_38_port, din(37) => 
                           state_main_in_p1_37_port, din(36) => 
                           state_main_in_p1_36_port, din(35) => 
                           state_main_in_p1_35_port, din(34) => 
                           state_main_in_p1_34_port, din(33) => 
                           state_main_in_p1_33_port, din(32) => 
                           state_main_in_p1_32_port, din(31) => 
                           state_main_in_p1_31_port, din(30) => 
                           state_main_in_p1_30_port, din(29) => 
                           state_main_in_p1_29_port, din(28) => 
                           state_main_in_p1_28_port, din(27) => 
                           state_main_in_p1_27_port, din(26) => 
                           state_main_in_p1_26_port, din(25) => 
                           state_main_in_p1_25_port, din(24) => 
                           state_main_in_p1_24_port, din(23) => 
                           state_main_in_p1_23_port, din(22) => 
                           state_main_in_p1_22_port, din(21) => 
                           state_main_in_p1_21_port, din(20) => 
                           state_main_in_p1_20_port, din(19) => 
                           state_main_in_p1_19_port, din(18) => 
                           state_main_in_p1_18_port, din(17) => 
                           state_main_in_p1_17_port, din(16) => 
                           state_main_in_p1_16_port, din(15) => 
                           state_main_in_p1_15_port, din(14) => 
                           state_main_in_p1_14_port, din(13) => 
                           state_main_in_p1_13_port, din(12) => 
                           state_main_in_p1_12_port, din(11) => 
                           state_main_in_p1_11_port, din(10) => 
                           state_main_in_p1_10_port, din(9) => 
                           state_main_in_p1_9_port, din(8) => 
                           state_main_in_p1_8_port, din(7) => 
                           state_main_in_p1_7_port, din(6) => 
                           state_main_in_p1_6_port, din(5) => 
                           state_main_in_p1_5_port, din(4) => 
                           state_main_in_p1_4_port, din(3) => 
                           state_main_in_p1_3_port, din(2) => 
                           state_main_in_p1_2_port, din(1) => 
                           state_main_in_p1_1_port, din(0) => 
                           state_main_in_p1_0_port, qout(127) => 
                           state_main_out_plane1_127_port, qout(126) => 
                           state_main_out_plane1_126_port, qout(125) => 
                           state_main_out_plane1_125_port, qout(124) => 
                           state_main_out_plane1_124_port, qout(123) => 
                           state_main_out_plane1_123_port, qout(122) => 
                           state_main_out_plane1_122_port, qout(121) => 
                           state_main_out_plane1_121_port, qout(120) => 
                           state_main_out_plane1_120_port, qout(119) => 
                           state_main_out_plane1_119_port, qout(118) => 
                           state_main_out_plane1_118_port, qout(117) => 
                           state_main_out_plane1_117_port, qout(116) => 
                           state_main_out_plane1_116_port, qout(115) => 
                           state_main_out_plane1_115_port, qout(114) => 
                           state_main_out_plane1_114_port, qout(113) => 
                           state_main_out_plane1_113_port, qout(112) => 
                           state_main_out_plane1_112_port, qout(111) => 
                           state_main_out_plane1_111_port, qout(110) => 
                           state_main_out_plane1_110_port, qout(109) => 
                           state_main_out_plane1_109_port, qout(108) => 
                           state_main_out_plane1_108_port, qout(107) => 
                           state_main_out_plane1_107_port, qout(106) => 
                           state_main_out_plane1_106_port, qout(105) => 
                           state_main_out_plane1_105_port, qout(104) => 
                           state_main_out_plane1_104_port, qout(103) => 
                           state_main_out_plane1_103_port, qout(102) => 
                           state_main_out_plane1_102_port, qout(101) => 
                           state_main_out_plane1_101_port, qout(100) => 
                           state_main_out_plane1_100_port, qout(99) => 
                           state_main_out_plane1_99_port, qout(98) => 
                           state_main_out_plane1_98_port, qout(97) => 
                           state_main_out_plane1_97_port, qout(96) => 
                           state_main_out_plane1_96_port, qout(95) => 
                           state_main_out_plane1_95_port, qout(94) => 
                           state_main_out_plane1_94_port, qout(93) => 
                           state_main_out_plane1_93_port, qout(92) => 
                           state_main_out_plane1_92_port, qout(91) => 
                           state_main_out_plane1_91_port, qout(90) => 
                           state_main_out_plane1_90_port, qout(89) => 
                           state_main_out_plane1_89_port, qout(88) => 
                           state_main_out_plane1_88_port, qout(87) => 
                           state_main_out_plane1_87_port, qout(86) => 
                           state_main_out_plane1_86_port, qout(85) => 
                           state_main_out_plane1_85_port, qout(84) => 
                           state_main_out_plane1_84_port, qout(83) => 
                           state_main_out_plane1_83_port, qout(82) => 
                           state_main_out_plane1_82_port, qout(81) => 
                           state_main_out_plane1_81_port, qout(80) => 
                           state_main_out_plane1_80_port, qout(79) => 
                           state_main_out_plane1_79_port, qout(78) => 
                           state_main_out_plane1_78_port, qout(77) => 
                           state_main_out_plane1_77_port, qout(76) => 
                           state_main_out_plane1_76_port, qout(75) => 
                           state_main_out_plane1_75_port, qout(74) => 
                           state_main_out_plane1_74_port, qout(73) => 
                           state_main_out_plane1_73_port, qout(72) => 
                           state_main_out_plane1_72_port, qout(71) => 
                           state_main_out_plane1_71_port, qout(70) => 
                           state_main_out_plane1_70_port, qout(69) => 
                           state_main_out_plane1_69_port, qout(68) => 
                           state_main_out_plane1_68_port, qout(67) => 
                           state_main_out_plane1_67_port, qout(66) => 
                           state_main_out_plane1_66_port, qout(65) => 
                           state_main_out_plane1_65_port, qout(64) => 
                           state_main_out_plane1_64_port, qout(63) => 
                           state_main_out_plane1_63_port, qout(62) => 
                           state_main_out_plane1_62_port, qout(61) => 
                           state_main_out_plane1_61_port, qout(60) => 
                           state_main_out_plane1_60_port, qout(59) => 
                           state_main_out_plane1_59_port, qout(58) => 
                           state_main_out_plane1_58_port, qout(57) => 
                           state_main_out_plane1_57_port, qout(56) => 
                           state_main_out_plane1_56_port, qout(55) => 
                           state_main_out_plane1_55_port, qout(54) => 
                           state_main_out_plane1_54_port, qout(53) => 
                           state_main_out_plane1_53_port, qout(52) => 
                           state_main_out_plane1_52_port, qout(51) => 
                           state_main_out_plane1_51_port, qout(50) => 
                           state_main_out_plane1_50_port, qout(49) => 
                           state_main_out_plane1_49_port, qout(48) => 
                           state_main_out_plane1_48_port, qout(47) => 
                           state_main_out_plane1_47_port, qout(46) => 
                           state_main_out_plane1_46_port, qout(45) => 
                           state_main_out_plane1_45_port, qout(44) => 
                           state_main_out_plane1_44_port, qout(43) => 
                           state_main_out_plane1_43_port, qout(42) => 
                           state_main_out_plane1_42_port, qout(41) => 
                           state_main_out_plane1_41_port, qout(40) => 
                           state_main_out_plane1_40_port, qout(39) => 
                           state_main_out_plane1_39_port, qout(38) => 
                           state_main_out_plane1_38_port, qout(37) => 
                           state_main_out_plane1_37_port, qout(36) => 
                           state_main_out_plane1_36_port, qout(35) => 
                           state_main_out_plane1_35_port, qout(34) => 
                           state_main_out_plane1_34_port, qout(33) => 
                           state_main_out_plane1_33_port, qout(32) => 
                           state_main_out_plane1_32_port, qout(31) => 
                           state_main_out_plane1_31_port, qout(30) => 
                           state_main_out_plane1_30_port, qout(29) => 
                           state_main_out_plane1_29_port, qout(28) => 
                           state_main_out_plane1_28_port, qout(27) => 
                           state_main_out_plane1_27_port, qout(26) => 
                           state_main_out_plane1_26_port, qout(25) => 
                           state_main_out_plane1_25_port, qout(24) => 
                           state_main_out_plane1_24_port, qout(23) => 
                           state_main_out_plane1_23_port, qout(22) => 
                           state_main_out_plane1_22_port, qout(21) => 
                           state_main_out_plane1_21_port, qout(20) => 
                           state_main_out_plane1_20_port, qout(19) => 
                           state_main_out_plane1_19_port, qout(18) => 
                           state_main_out_plane1_18_port, qout(17) => 
                           state_main_out_plane1_17_port, qout(16) => 
                           state_main_out_plane1_16_port, qout(15) => 
                           state_main_out_plane1_15_port, qout(14) => 
                           state_main_out_plane1_14_port, qout(13) => 
                           state_main_out_plane1_13_port, qout(12) => 
                           state_main_out_plane1_12_port, qout(11) => 
                           state_main_out_plane1_11_port, qout(10) => 
                           state_main_out_plane1_10_port, qout(9) => 
                           state_main_out_plane1_9_port, qout(8) => 
                           state_main_out_plane1_8_port, qout(7) => 
                           state_main_out_plane1_7_port, qout(6) => 
                           state_main_out_plane1_6_port, qout(5) => 
                           state_main_out_plane1_5_port, qout(4) => 
                           state_main_out_plane1_4_port, qout(3) => 
                           state_main_out_plane1_3_port, qout(2) => 
                           state_main_out_plane1_2_port, qout(1) => 
                           state_main_out_plane1_1_port, qout(0) => 
                           state_main_out_plane1_0_port);
   state_main_p2 : reg_custom_LEN128_1 port map( clk => clk, en => 
                           state_main_en(2), din(127) => 
                           state_main_in_p2_127_port, din(126) => 
                           state_main_in_p2_126_port, din(125) => 
                           state_main_in_p2_125_port, din(124) => 
                           state_main_in_p2_124_port, din(123) => 
                           state_main_in_p2_123_port, din(122) => 
                           state_main_in_p2_122_port, din(121) => 
                           state_main_in_p2_121_port, din(120) => 
                           state_main_in_p2_120_port, din(119) => 
                           state_main_in_p2_119_port, din(118) => 
                           state_main_in_p2_118_port, din(117) => 
                           state_main_in_p2_117_port, din(116) => 
                           state_main_in_p2_116_port, din(115) => 
                           state_main_in_p2_115_port, din(114) => 
                           state_main_in_p2_114_port, din(113) => 
                           state_main_in_p2_113_port, din(112) => 
                           state_main_in_p2_112_port, din(111) => 
                           state_main_in_p2_111_port, din(110) => 
                           state_main_in_p2_110_port, din(109) => 
                           state_main_in_p2_109_port, din(108) => 
                           state_main_in_p2_108_port, din(107) => 
                           state_main_in_p2_107_port, din(106) => 
                           state_main_in_p2_106_port, din(105) => 
                           state_main_in_p2_105_port, din(104) => 
                           state_main_in_p2_104_port, din(103) => 
                           state_main_in_p2_103_port, din(102) => 
                           state_main_in_p2_102_port, din(101) => 
                           state_main_in_p2_101_port, din(100) => 
                           state_main_in_p2_100_port, din(99) => 
                           state_main_in_p2_99_port, din(98) => 
                           state_main_in_p2_98_port, din(97) => 
                           state_main_in_p2_97_port, din(96) => 
                           state_main_in_p2_96_port, din(95) => 
                           state_main_in_p2_95_port, din(94) => 
                           state_main_in_p2_94_port, din(93) => 
                           state_main_in_p2_93_port, din(92) => 
                           state_main_in_p2_92_port, din(91) => 
                           state_main_in_p2_91_port, din(90) => 
                           state_main_in_p2_90_port, din(89) => 
                           state_main_in_p2_89_port, din(88) => 
                           state_main_in_p2_88_port, din(87) => 
                           state_main_in_p2_87_port, din(86) => 
                           state_main_in_p2_86_port, din(85) => 
                           state_main_in_p2_85_port, din(84) => 
                           state_main_in_p2_84_port, din(83) => 
                           state_main_in_p2_83_port, din(82) => 
                           state_main_in_p2_82_port, din(81) => 
                           state_main_in_p2_81_port, din(80) => 
                           state_main_in_p2_80_port, din(79) => 
                           state_main_in_p2_79_port, din(78) => 
                           state_main_in_p2_78_port, din(77) => 
                           state_main_in_p2_77_port, din(76) => 
                           state_main_in_p2_76_port, din(75) => 
                           state_main_in_p2_75_port, din(74) => 
                           state_main_in_p2_74_port, din(73) => 
                           state_main_in_p2_73_port, din(72) => 
                           state_main_in_p2_72_port, din(71) => 
                           state_main_in_p2_71_port, din(70) => 
                           state_main_in_p2_70_port, din(69) => 
                           state_main_in_p2_69_port, din(68) => 
                           state_main_in_p2_68_port, din(67) => 
                           state_main_in_p2_67_port, din(66) => 
                           state_main_in_p2_66_port, din(65) => 
                           state_main_in_p2_65_port, din(64) => 
                           state_main_in_p2_64_port, din(63) => 
                           state_main_in_p2_63_port, din(62) => 
                           state_main_in_p2_62_port, din(61) => 
                           state_main_in_p2_61_port, din(60) => 
                           state_main_in_p2_60_port, din(59) => 
                           state_main_in_p2_59_port, din(58) => 
                           state_main_in_p2_58_port, din(57) => 
                           state_main_in_p2_57_port, din(56) => 
                           state_main_in_p2_56_port, din(55) => 
                           state_main_in_p2_55_port, din(54) => 
                           state_main_in_p2_54_port, din(53) => 
                           state_main_in_p2_53_port, din(52) => 
                           state_main_in_p2_52_port, din(51) => 
                           state_main_in_p2_51_port, din(50) => 
                           state_main_in_p2_50_port, din(49) => 
                           state_main_in_p2_49_port, din(48) => 
                           state_main_in_p2_48_port, din(47) => 
                           state_main_in_p2_47_port, din(46) => 
                           state_main_in_p2_46_port, din(45) => 
                           state_main_in_p2_45_port, din(44) => 
                           state_main_in_p2_44_port, din(43) => 
                           state_main_in_p2_43_port, din(42) => 
                           state_main_in_p2_42_port, din(41) => 
                           state_main_in_p2_41_port, din(40) => 
                           state_main_in_p2_40_port, din(39) => 
                           state_main_in_p2_39_port, din(38) => 
                           state_main_in_p2_38_port, din(37) => 
                           state_main_in_p2_37_port, din(36) => 
                           state_main_in_p2_36_port, din(35) => 
                           state_main_in_p2_35_port, din(34) => 
                           state_main_in_p2_34_port, din(33) => 
                           state_main_in_p2_33_port, din(32) => 
                           state_main_in_p2_32_port, din(31) => 
                           state_main_in_p2_31_port, din(30) => 
                           state_main_in_p2_30_port, din(29) => 
                           state_main_in_p2_29_port, din(28) => 
                           state_main_in_p2_28_port, din(27) => 
                           state_main_in_p2_27_port, din(26) => 
                           state_main_in_p2_26_port, din(25) => 
                           state_main_in_p2_25_port, din(24) => 
                           state_main_in_p2_24_port, din(23) => 
                           state_main_in_p2_23_port, din(22) => 
                           state_main_in_p2_22_port, din(21) => 
                           state_main_in_p2_21_port, din(20) => 
                           state_main_in_p2_20_port, din(19) => 
                           state_main_in_p2_19_port, din(18) => 
                           state_main_in_p2_18_port, din(17) => 
                           state_main_in_p2_17_port, din(16) => 
                           state_main_in_p2_16_port, din(15) => 
                           state_main_in_p2_15_port, din(14) => 
                           state_main_in_p2_14_port, din(13) => 
                           state_main_in_p2_13_port, din(12) => 
                           state_main_in_p2_12_port, din(11) => 
                           state_main_in_p2_11_port, din(10) => 
                           state_main_in_p2_10_port, din(9) => 
                           state_main_in_p2_9_port, din(8) => 
                           state_main_in_p2_8_port, din(7) => 
                           state_main_in_p2_7_port, din(6) => 
                           state_main_in_p2_6_port, din(5) => 
                           state_main_in_p2_5_port, din(4) => 
                           state_main_in_p2_4_port, din(3) => 
                           state_main_in_p2_3_port, din(2) => 
                           state_main_in_p2_2_port, din(1) => 
                           state_main_in_p2_1_port, din(0) => 
                           state_main_in_p2_0_port, qout(127) => 
                           state_main_out_plane2_127_port, qout(126) => 
                           state_main_out_plane2_126_port, qout(125) => 
                           state_main_out_plane2_125_port, qout(124) => 
                           state_main_out_plane2_124_port, qout(123) => 
                           state_main_out_plane2_123_port, qout(122) => 
                           state_main_out_plane2_122_port, qout(121) => 
                           state_main_out_plane2_121_port, qout(120) => 
                           state_main_out_plane2_120_port, qout(119) => 
                           state_main_out_plane2_119_port, qout(118) => 
                           state_main_out_plane2_118_port, qout(117) => 
                           state_main_out_plane2_117_port, qout(116) => 
                           state_main_out_plane2_116_port, qout(115) => 
                           state_main_out_plane2_115_port, qout(114) => 
                           state_main_out_plane2_114_port, qout(113) => 
                           state_main_out_plane2_113_port, qout(112) => 
                           state_main_out_plane2_112_port, qout(111) => 
                           state_main_out_plane2_111_port, qout(110) => 
                           state_main_out_plane2_110_port, qout(109) => 
                           state_main_out_plane2_109_port, qout(108) => 
                           state_main_out_plane2_108_port, qout(107) => 
                           state_main_out_plane2_107_port, qout(106) => 
                           state_main_out_plane2_106_port, qout(105) => 
                           state_main_out_plane2_105_port, qout(104) => 
                           state_main_out_plane2_104_port, qout(103) => 
                           state_main_out_plane2_103_port, qout(102) => 
                           state_main_out_plane2_102_port, qout(101) => 
                           state_main_out_plane2_101_port, qout(100) => 
                           state_main_out_plane2_100_port, qout(99) => 
                           state_main_out_plane2_99_port, qout(98) => 
                           state_main_out_plane2_98_port, qout(97) => 
                           state_main_out_plane2_97_port, qout(96) => 
                           state_main_out_plane2_96_port, qout(95) => 
                           state_main_out_plane2_95_port, qout(94) => 
                           state_main_out_plane2_94_port, qout(93) => 
                           state_main_out_plane2_93_port, qout(92) => 
                           state_main_out_plane2_92_port, qout(91) => 
                           state_main_out_plane2_91_port, qout(90) => 
                           state_main_out_plane2_90_port, qout(89) => 
                           state_main_out_plane2_89_port, qout(88) => 
                           state_main_out_plane2_88_port, qout(87) => 
                           state_main_out_plane2_87_port, qout(86) => 
                           state_main_out_plane2_86_port, qout(85) => 
                           state_main_out_plane2_85_port, qout(84) => 
                           state_main_out_plane2_84_port, qout(83) => 
                           state_main_out_plane2_83_port, qout(82) => 
                           state_main_out_plane2_82_port, qout(81) => 
                           state_main_out_plane2_81_port, qout(80) => 
                           state_main_out_plane2_80_port, qout(79) => 
                           state_main_out_plane2_79_port, qout(78) => 
                           state_main_out_plane2_78_port, qout(77) => 
                           state_main_out_plane2_77_port, qout(76) => 
                           state_main_out_plane2_76_port, qout(75) => 
                           state_main_out_plane2_75_port, qout(74) => 
                           state_main_out_plane2_74_port, qout(73) => 
                           state_main_out_plane2_73_port, qout(72) => 
                           state_main_out_plane2_72_port, qout(71) => 
                           state_main_out_plane2_71_port, qout(70) => 
                           state_main_out_plane2_70_port, qout(69) => 
                           state_main_out_plane2_69_port, qout(68) => 
                           state_main_out_plane2_68_port, qout(67) => 
                           state_main_out_plane2_67_port, qout(66) => 
                           state_main_out_plane2_66_port, qout(65) => 
                           state_main_out_plane2_65_port, qout(64) => 
                           state_main_out_plane2_64_port, qout(63) => 
                           state_main_out_plane2_63_port, qout(62) => 
                           state_main_out_plane2_62_port, qout(61) => 
                           state_main_out_plane2_61_port, qout(60) => 
                           state_main_out_plane2_60_port, qout(59) => 
                           state_main_out_plane2_59_port, qout(58) => 
                           state_main_out_plane2_58_port, qout(57) => 
                           state_main_out_plane2_57_port, qout(56) => 
                           state_main_out_plane2_56_port, qout(55) => 
                           state_main_out_plane2_55_port, qout(54) => 
                           state_main_out_plane2_54_port, qout(53) => 
                           state_main_out_plane2_53_port, qout(52) => 
                           state_main_out_plane2_52_port, qout(51) => 
                           state_main_out_plane2_51_port, qout(50) => 
                           state_main_out_plane2_50_port, qout(49) => 
                           state_main_out_plane2_49_port, qout(48) => 
                           state_main_out_plane2_48_port, qout(47) => 
                           state_main_out_plane2_47_port, qout(46) => 
                           state_main_out_plane2_46_port, qout(45) => 
                           state_main_out_plane2_45_port, qout(44) => 
                           state_main_out_plane2_44_port, qout(43) => 
                           state_main_out_plane2_43_port, qout(42) => 
                           state_main_out_plane2_42_port, qout(41) => 
                           state_main_out_plane2_41_port, qout(40) => 
                           state_main_out_plane2_40_port, qout(39) => 
                           state_main_out_plane2_39_port, qout(38) => 
                           state_main_out_plane2_38_port, qout(37) => 
                           state_main_out_plane2_37_port, qout(36) => 
                           state_main_out_plane2_36_port, qout(35) => 
                           state_main_out_plane2_35_port, qout(34) => 
                           state_main_out_plane2_34_port, qout(33) => 
                           state_main_out_plane2_33_port, qout(32) => 
                           state_main_out_plane2_32_port, qout(31) => 
                           state_main_out_plane2_31_port, qout(30) => 
                           state_main_out_plane2_30_port, qout(29) => 
                           state_main_out_plane2_29_port, qout(28) => 
                           state_main_out_plane2_28_port, qout(27) => 
                           state_main_out_plane2_27_port, qout(26) => 
                           state_main_out_plane2_26_port, qout(25) => 
                           state_main_out_plane2_25_port, qout(24) => 
                           state_main_out_plane2_24_port, qout(23) => 
                           state_main_out_plane2_23_port, qout(22) => 
                           state_main_out_plane2_22_port, qout(21) => 
                           state_main_out_plane2_21_port, qout(20) => 
                           state_main_out_plane2_20_port, qout(19) => 
                           state_main_out_plane2_19_port, qout(18) => 
                           state_main_out_plane2_18_port, qout(17) => 
                           state_main_out_plane2_17_port, qout(16) => 
                           state_main_out_plane2_16_port, qout(15) => 
                           state_main_out_plane2_15_port, qout(14) => 
                           state_main_out_plane2_14_port, qout(13) => 
                           state_main_out_plane2_13_port, qout(12) => 
                           state_main_out_plane2_12_port, qout(11) => 
                           state_main_out_plane2_11_port, qout(10) => 
                           state_main_out_plane2_10_port, qout(9) => 
                           state_main_out_plane2_9_port, qout(8) => 
                           state_main_out_plane2_8_port, qout(7) => 
                           state_main_out_plane2_7_port, qout(6) => 
                           state_main_out_plane2_6_port, qout(5) => 
                           state_main_out_plane2_5_port, qout(4) => 
                           state_main_out_plane2_4_port, qout(3) => 
                           state_main_out_plane2_3_port, qout(2) => 
                           state_main_out_plane2_2_port, qout(1) => 
                           state_main_out_plane2_1_port, qout(0) => 
                           state_main_out_plane2_0_port);
   XOODOO_PERM : xoodoo_round_ADDRESS_LEN384_1 port map( INPUT(383) => 
                           state_main_out_plane2_127_port, INPUT(382) => 
                           state_main_out_plane2_126_port, INPUT(381) => 
                           state_main_out_plane2_125_port, INPUT(380) => 
                           state_main_out_plane2_124_port, INPUT(379) => 
                           state_main_out_plane2_123_port, INPUT(378) => 
                           state_main_out_plane2_122_port, INPUT(377) => 
                           state_main_out_plane2_121_port, INPUT(376) => 
                           state_main_out_plane2_120_port, INPUT(375) => 
                           state_main_out_plane2_119_port, INPUT(374) => 
                           state_main_out_plane2_118_port, INPUT(373) => 
                           state_main_out_plane2_117_port, INPUT(372) => 
                           state_main_out_plane2_116_port, INPUT(371) => 
                           state_main_out_plane2_115_port, INPUT(370) => 
                           state_main_out_plane2_114_port, INPUT(369) => 
                           state_main_out_plane2_113_port, INPUT(368) => 
                           state_main_out_plane2_112_port, INPUT(367) => 
                           state_main_out_plane2_111_port, INPUT(366) => 
                           state_main_out_plane2_110_port, INPUT(365) => 
                           state_main_out_plane2_109_port, INPUT(364) => 
                           state_main_out_plane2_108_port, INPUT(363) => 
                           state_main_out_plane2_107_port, INPUT(362) => 
                           state_main_out_plane2_106_port, INPUT(361) => 
                           state_main_out_plane2_105_port, INPUT(360) => 
                           state_main_out_plane2_104_port, INPUT(359) => 
                           state_main_out_plane2_103_port, INPUT(358) => 
                           state_main_out_plane2_102_port, INPUT(357) => 
                           state_main_out_plane2_101_port, INPUT(356) => 
                           state_main_out_plane2_100_port, INPUT(355) => 
                           state_main_out_plane2_99_port, INPUT(354) => 
                           state_main_out_plane2_98_port, INPUT(353) => 
                           state_main_out_plane2_97_port, INPUT(352) => 
                           state_main_out_plane2_96_port, INPUT(351) => 
                           state_main_out_plane2_95_port, INPUT(350) => 
                           state_main_out_plane2_94_port, INPUT(349) => 
                           state_main_out_plane2_93_port, INPUT(348) => 
                           state_main_out_plane2_92_port, INPUT(347) => 
                           state_main_out_plane2_91_port, INPUT(346) => 
                           state_main_out_plane2_90_port, INPUT(345) => 
                           state_main_out_plane2_89_port, INPUT(344) => 
                           state_main_out_plane2_88_port, INPUT(343) => 
                           state_main_out_plane2_87_port, INPUT(342) => 
                           state_main_out_plane2_86_port, INPUT(341) => 
                           state_main_out_plane2_85_port, INPUT(340) => 
                           state_main_out_plane2_84_port, INPUT(339) => 
                           state_main_out_plane2_83_port, INPUT(338) => 
                           state_main_out_plane2_82_port, INPUT(337) => 
                           state_main_out_plane2_81_port, INPUT(336) => 
                           state_main_out_plane2_80_port, INPUT(335) => 
                           state_main_out_plane2_79_port, INPUT(334) => 
                           state_main_out_plane2_78_port, INPUT(333) => 
                           state_main_out_plane2_77_port, INPUT(332) => 
                           state_main_out_plane2_76_port, INPUT(331) => 
                           state_main_out_plane2_75_port, INPUT(330) => 
                           state_main_out_plane2_74_port, INPUT(329) => 
                           state_main_out_plane2_73_port, INPUT(328) => 
                           state_main_out_plane2_72_port, INPUT(327) => 
                           state_main_out_plane2_71_port, INPUT(326) => 
                           state_main_out_plane2_70_port, INPUT(325) => 
                           state_main_out_plane2_69_port, INPUT(324) => 
                           state_main_out_plane2_68_port, INPUT(323) => 
                           state_main_out_plane2_67_port, INPUT(322) => 
                           state_main_out_plane2_66_port, INPUT(321) => 
                           state_main_out_plane2_65_port, INPUT(320) => 
                           state_main_out_plane2_64_port, INPUT(319) => 
                           state_main_out_plane2_63_port, INPUT(318) => 
                           state_main_out_plane2_62_port, INPUT(317) => 
                           state_main_out_plane2_61_port, INPUT(316) => 
                           state_main_out_plane2_60_port, INPUT(315) => 
                           state_main_out_plane2_59_port, INPUT(314) => 
                           state_main_out_plane2_58_port, INPUT(313) => 
                           state_main_out_plane2_57_port, INPUT(312) => 
                           state_main_out_plane2_56_port, INPUT(311) => 
                           state_main_out_plane2_55_port, INPUT(310) => 
                           state_main_out_plane2_54_port, INPUT(309) => 
                           state_main_out_plane2_53_port, INPUT(308) => 
                           state_main_out_plane2_52_port, INPUT(307) => 
                           state_main_out_plane2_51_port, INPUT(306) => 
                           state_main_out_plane2_50_port, INPUT(305) => 
                           state_main_out_plane2_49_port, INPUT(304) => 
                           state_main_out_plane2_48_port, INPUT(303) => 
                           state_main_out_plane2_47_port, INPUT(302) => 
                           state_main_out_plane2_46_port, INPUT(301) => 
                           state_main_out_plane2_45_port, INPUT(300) => 
                           state_main_out_plane2_44_port, INPUT(299) => 
                           state_main_out_plane2_43_port, INPUT(298) => 
                           state_main_out_plane2_42_port, INPUT(297) => 
                           state_main_out_plane2_41_port, INPUT(296) => 
                           state_main_out_plane2_40_port, INPUT(295) => 
                           state_main_out_plane2_39_port, INPUT(294) => 
                           state_main_out_plane2_38_port, INPUT(293) => 
                           state_main_out_plane2_37_port, INPUT(292) => 
                           state_main_out_plane2_36_port, INPUT(291) => 
                           state_main_out_plane2_35_port, INPUT(290) => 
                           state_main_out_plane2_34_port, INPUT(289) => 
                           state_main_out_plane2_33_port, INPUT(288) => 
                           state_main_out_plane2_32_port, INPUT(287) => 
                           state_main_out_plane2_31_port, INPUT(286) => 
                           state_main_out_plane2_30_port, INPUT(285) => 
                           state_main_out_plane2_29_port, INPUT(284) => 
                           state_main_out_plane2_28_port, INPUT(283) => 
                           state_main_out_plane2_27_port, INPUT(282) => 
                           state_main_out_plane2_26_port, INPUT(281) => 
                           state_main_out_plane2_25_port, INPUT(280) => 
                           state_main_out_plane2_24_port, INPUT(279) => 
                           state_main_out_plane2_23_port, INPUT(278) => 
                           state_main_out_plane2_22_port, INPUT(277) => 
                           state_main_out_plane2_21_port, INPUT(276) => 
                           state_main_out_plane2_20_port, INPUT(275) => 
                           state_main_out_plane2_19_port, INPUT(274) => 
                           state_main_out_plane2_18_port, INPUT(273) => 
                           state_main_out_plane2_17_port, INPUT(272) => 
                           state_main_out_plane2_16_port, INPUT(271) => 
                           state_main_out_plane2_15_port, INPUT(270) => 
                           state_main_out_plane2_14_port, INPUT(269) => 
                           state_main_out_plane2_13_port, INPUT(268) => 
                           state_main_out_plane2_12_port, INPUT(267) => 
                           state_main_out_plane2_11_port, INPUT(266) => 
                           state_main_out_plane2_10_port, INPUT(265) => 
                           state_main_out_plane2_9_port, INPUT(264) => 
                           state_main_out_plane2_8_port, INPUT(263) => 
                           state_main_out_plane2_7_port, INPUT(262) => 
                           state_main_out_plane2_6_port, INPUT(261) => 
                           state_main_out_plane2_5_port, INPUT(260) => 
                           state_main_out_plane2_4_port, INPUT(259) => 
                           state_main_out_plane2_3_port, INPUT(258) => 
                           state_main_out_plane2_2_port, INPUT(257) => 
                           state_main_out_plane2_1_port, INPUT(256) => 
                           state_main_out_plane2_0_port, INPUT(255) => 
                           state_main_out_plane1_127_port, INPUT(254) => 
                           state_main_out_plane1_126_port, INPUT(253) => 
                           state_main_out_plane1_125_port, INPUT(252) => 
                           state_main_out_plane1_124_port, INPUT(251) => 
                           state_main_out_plane1_123_port, INPUT(250) => 
                           state_main_out_plane1_122_port, INPUT(249) => 
                           state_main_out_plane1_121_port, INPUT(248) => 
                           state_main_out_plane1_120_port, INPUT(247) => 
                           state_main_out_plane1_119_port, INPUT(246) => 
                           state_main_out_plane1_118_port, INPUT(245) => 
                           state_main_out_plane1_117_port, INPUT(244) => 
                           state_main_out_plane1_116_port, INPUT(243) => 
                           state_main_out_plane1_115_port, INPUT(242) => 
                           state_main_out_plane1_114_port, INPUT(241) => 
                           state_main_out_plane1_113_port, INPUT(240) => 
                           state_main_out_plane1_112_port, INPUT(239) => 
                           state_main_out_plane1_111_port, INPUT(238) => 
                           state_main_out_plane1_110_port, INPUT(237) => 
                           state_main_out_plane1_109_port, INPUT(236) => 
                           state_main_out_plane1_108_port, INPUT(235) => 
                           state_main_out_plane1_107_port, INPUT(234) => 
                           state_main_out_plane1_106_port, INPUT(233) => 
                           state_main_out_plane1_105_port, INPUT(232) => 
                           state_main_out_plane1_104_port, INPUT(231) => 
                           state_main_out_plane1_103_port, INPUT(230) => 
                           state_main_out_plane1_102_port, INPUT(229) => 
                           state_main_out_plane1_101_port, INPUT(228) => 
                           state_main_out_plane1_100_port, INPUT(227) => 
                           state_main_out_plane1_99_port, INPUT(226) => 
                           state_main_out_plane1_98_port, INPUT(225) => 
                           state_main_out_plane1_97_port, INPUT(224) => 
                           state_main_out_plane1_96_port, INPUT(223) => 
                           state_main_out_plane1_95_port, INPUT(222) => 
                           state_main_out_plane1_94_port, INPUT(221) => 
                           state_main_out_plane1_93_port, INPUT(220) => 
                           state_main_out_plane1_92_port, INPUT(219) => 
                           state_main_out_plane1_91_port, INPUT(218) => 
                           state_main_out_plane1_90_port, INPUT(217) => 
                           state_main_out_plane1_89_port, INPUT(216) => 
                           state_main_out_plane1_88_port, INPUT(215) => 
                           state_main_out_plane1_87_port, INPUT(214) => 
                           state_main_out_plane1_86_port, INPUT(213) => 
                           state_main_out_plane1_85_port, INPUT(212) => 
                           state_main_out_plane1_84_port, INPUT(211) => 
                           state_main_out_plane1_83_port, INPUT(210) => 
                           state_main_out_plane1_82_port, INPUT(209) => 
                           state_main_out_plane1_81_port, INPUT(208) => 
                           state_main_out_plane1_80_port, INPUT(207) => 
                           state_main_out_plane1_79_port, INPUT(206) => 
                           state_main_out_plane1_78_port, INPUT(205) => 
                           state_main_out_plane1_77_port, INPUT(204) => 
                           state_main_out_plane1_76_port, INPUT(203) => 
                           state_main_out_plane1_75_port, INPUT(202) => 
                           state_main_out_plane1_74_port, INPUT(201) => 
                           state_main_out_plane1_73_port, INPUT(200) => 
                           state_main_out_plane1_72_port, INPUT(199) => 
                           state_main_out_plane1_71_port, INPUT(198) => 
                           state_main_out_plane1_70_port, INPUT(197) => 
                           state_main_out_plane1_69_port, INPUT(196) => 
                           state_main_out_plane1_68_port, INPUT(195) => 
                           state_main_out_plane1_67_port, INPUT(194) => 
                           state_main_out_plane1_66_port, INPUT(193) => 
                           state_main_out_plane1_65_port, INPUT(192) => 
                           state_main_out_plane1_64_port, INPUT(191) => 
                           state_main_out_plane1_63_port, INPUT(190) => 
                           state_main_out_plane1_62_port, INPUT(189) => 
                           state_main_out_plane1_61_port, INPUT(188) => 
                           state_main_out_plane1_60_port, INPUT(187) => 
                           state_main_out_plane1_59_port, INPUT(186) => 
                           state_main_out_plane1_58_port, INPUT(185) => 
                           state_main_out_plane1_57_port, INPUT(184) => 
                           state_main_out_plane1_56_port, INPUT(183) => 
                           state_main_out_plane1_55_port, INPUT(182) => 
                           state_main_out_plane1_54_port, INPUT(181) => 
                           state_main_out_plane1_53_port, INPUT(180) => 
                           state_main_out_plane1_52_port, INPUT(179) => 
                           state_main_out_plane1_51_port, INPUT(178) => 
                           state_main_out_plane1_50_port, INPUT(177) => 
                           state_main_out_plane1_49_port, INPUT(176) => 
                           state_main_out_plane1_48_port, INPUT(175) => 
                           state_main_out_plane1_47_port, INPUT(174) => 
                           state_main_out_plane1_46_port, INPUT(173) => 
                           state_main_out_plane1_45_port, INPUT(172) => 
                           state_main_out_plane1_44_port, INPUT(171) => 
                           state_main_out_plane1_43_port, INPUT(170) => 
                           state_main_out_plane1_42_port, INPUT(169) => 
                           state_main_out_plane1_41_port, INPUT(168) => 
                           state_main_out_plane1_40_port, INPUT(167) => 
                           state_main_out_plane1_39_port, INPUT(166) => 
                           state_main_out_plane1_38_port, INPUT(165) => 
                           state_main_out_plane1_37_port, INPUT(164) => 
                           state_main_out_plane1_36_port, INPUT(163) => 
                           state_main_out_plane1_35_port, INPUT(162) => 
                           state_main_out_plane1_34_port, INPUT(161) => 
                           state_main_out_plane1_33_port, INPUT(160) => 
                           state_main_out_plane1_32_port, INPUT(159) => 
                           state_main_out_plane1_31_port, INPUT(158) => 
                           state_main_out_plane1_30_port, INPUT(157) => 
                           state_main_out_plane1_29_port, INPUT(156) => 
                           state_main_out_plane1_28_port, INPUT(155) => 
                           state_main_out_plane1_27_port, INPUT(154) => 
                           state_main_out_plane1_26_port, INPUT(153) => 
                           state_main_out_plane1_25_port, INPUT(152) => 
                           state_main_out_plane1_24_port, INPUT(151) => 
                           state_main_out_plane1_23_port, INPUT(150) => 
                           state_main_out_plane1_22_port, INPUT(149) => 
                           state_main_out_plane1_21_port, INPUT(148) => 
                           state_main_out_plane1_20_port, INPUT(147) => 
                           state_main_out_plane1_19_port, INPUT(146) => 
                           state_main_out_plane1_18_port, INPUT(145) => 
                           state_main_out_plane1_17_port, INPUT(144) => 
                           state_main_out_plane1_16_port, INPUT(143) => 
                           state_main_out_plane1_15_port, INPUT(142) => 
                           state_main_out_plane1_14_port, INPUT(141) => 
                           state_main_out_plane1_13_port, INPUT(140) => 
                           state_main_out_plane1_12_port, INPUT(139) => 
                           state_main_out_plane1_11_port, INPUT(138) => 
                           state_main_out_plane1_10_port, INPUT(137) => 
                           state_main_out_plane1_9_port, INPUT(136) => 
                           state_main_out_plane1_8_port, INPUT(135) => 
                           state_main_out_plane1_7_port, INPUT(134) => 
                           state_main_out_plane1_6_port, INPUT(133) => 
                           state_main_out_plane1_5_port, INPUT(132) => 
                           state_main_out_plane1_4_port, INPUT(131) => 
                           state_main_out_plane1_3_port, INPUT(130) => 
                           state_main_out_plane1_2_port, INPUT(129) => 
                           state_main_out_plane1_1_port, INPUT(128) => 
                           state_main_out_plane1_0_port, INPUT(127) => 
                           state_main_out_plane0_127_port, INPUT(126) => 
                           state_main_out_plane0_126_port, INPUT(125) => 
                           state_main_out_plane0_125_port, INPUT(124) => 
                           state_main_out_plane0_124_port, INPUT(123) => 
                           state_main_out_plane0_123_port, INPUT(122) => 
                           state_main_out_plane0_122_port, INPUT(121) => 
                           state_main_out_plane0_121_port, INPUT(120) => 
                           state_main_out_plane0_120_port, INPUT(119) => 
                           state_main_out_plane0_119_port, INPUT(118) => 
                           state_main_out_plane0_118_port, INPUT(117) => 
                           state_main_out_plane0_117_port, INPUT(116) => 
                           state_main_out_plane0_116_port, INPUT(115) => 
                           state_main_out_plane0_115_port, INPUT(114) => 
                           state_main_out_plane0_114_port, INPUT(113) => 
                           state_main_out_plane0_113_port, INPUT(112) => 
                           state_main_out_plane0_112_port, INPUT(111) => 
                           state_main_out_plane0_111_port, INPUT(110) => 
                           state_main_out_plane0_110_port, INPUT(109) => 
                           state_main_out_plane0_109_port, INPUT(108) => 
                           state_main_out_plane0_108_port, INPUT(107) => 
                           state_main_out_plane0_107_port, INPUT(106) => 
                           state_main_out_plane0_106_port, INPUT(105) => 
                           state_main_out_plane0_105_port, INPUT(104) => 
                           state_main_out_plane0_104_port, INPUT(103) => 
                           state_main_out_plane0_103_port, INPUT(102) => 
                           state_main_out_plane0_102_port, INPUT(101) => 
                           state_main_out_plane0_101_port, INPUT(100) => 
                           state_main_out_plane0_100_port, INPUT(99) => 
                           state_main_out_plane0_99_port, INPUT(98) => 
                           state_main_out_plane0_98_port, INPUT(97) => 
                           state_main_out_plane0_97_port, INPUT(96) => 
                           state_main_out_plane0_96_port, INPUT(95) => 
                           state_main_out_plane0_95_port, INPUT(94) => 
                           state_main_out_plane0_94_port, INPUT(93) => 
                           state_main_out_plane0_93_port, INPUT(92) => 
                           state_main_out_plane0_92_port, INPUT(91) => 
                           state_main_out_plane0_91_port, INPUT(90) => 
                           state_main_out_plane0_90_port, INPUT(89) => 
                           state_main_out_plane0_89_port, INPUT(88) => 
                           state_main_out_plane0_88_port, INPUT(87) => 
                           state_main_out_plane0_87_port, INPUT(86) => 
                           state_main_out_plane0_86_port, INPUT(85) => 
                           state_main_out_plane0_85_port, INPUT(84) => 
                           state_main_out_plane0_84_port, INPUT(83) => 
                           state_main_out_plane0_83_port, INPUT(82) => 
                           state_main_out_plane0_82_port, INPUT(81) => 
                           state_main_out_plane0_81_port, INPUT(80) => 
                           state_main_out_plane0_80_port, INPUT(79) => 
                           state_main_out_plane0_79_port, INPUT(78) => 
                           state_main_out_plane0_78_port, INPUT(77) => 
                           state_main_out_plane0_77_port, INPUT(76) => 
                           state_main_out_plane0_76_port, INPUT(75) => 
                           state_main_out_plane0_75_port, INPUT(74) => 
                           state_main_out_plane0_74_port, INPUT(73) => 
                           state_main_out_plane0_73_port, INPUT(72) => 
                           state_main_out_plane0_72_port, INPUT(71) => 
                           state_main_out_plane0_71_port, INPUT(70) => 
                           state_main_out_plane0_70_port, INPUT(69) => 
                           state_main_out_plane0_69_port, INPUT(68) => 
                           state_main_out_plane0_68_port, INPUT(67) => 
                           state_main_out_plane0_67_port, INPUT(66) => 
                           state_main_out_plane0_66_port, INPUT(65) => 
                           state_main_out_plane0_65_port, INPUT(64) => 
                           state_main_out_plane0_64_port, INPUT(63) => 
                           state_main_out_plane0_63_port, INPUT(62) => 
                           state_main_out_plane0_62_port, INPUT(61) => 
                           state_main_out_plane0_61_port, INPUT(60) => 
                           state_main_out_plane0_60_port, INPUT(59) => 
                           state_main_out_plane0_59_port, INPUT(58) => 
                           state_main_out_plane0_58_port, INPUT(57) => 
                           state_main_out_plane0_57_port, INPUT(56) => 
                           state_main_out_plane0_56_port, INPUT(55) => 
                           state_main_out_plane0_55_port, INPUT(54) => 
                           state_main_out_plane0_54_port, INPUT(53) => 
                           state_main_out_plane0_53_port, INPUT(52) => 
                           state_main_out_plane0_52_port, INPUT(51) => 
                           state_main_out_plane0_51_port, INPUT(50) => 
                           state_main_out_plane0_50_port, INPUT(49) => 
                           state_main_out_plane0_49_port, INPUT(48) => 
                           state_main_out_plane0_48_port, INPUT(47) => 
                           state_main_out_plane0_47_port, INPUT(46) => 
                           state_main_out_plane0_46_port, INPUT(45) => 
                           state_main_out_plane0_45_port, INPUT(44) => 
                           state_main_out_plane0_44_port, INPUT(43) => 
                           state_main_out_plane0_43_port, INPUT(42) => 
                           state_main_out_plane0_42_port, INPUT(41) => 
                           state_main_out_plane0_41_port, INPUT(40) => 
                           state_main_out_plane0_40_port, INPUT(39) => 
                           state_main_out_plane0_39_port, INPUT(38) => 
                           state_main_out_plane0_38_port, INPUT(37) => 
                           state_main_out_plane0_37_port, INPUT(36) => 
                           state_main_out_plane0_36_port, INPUT(35) => 
                           state_main_out_plane0_35_port, INPUT(34) => 
                           state_main_out_plane0_34_port, INPUT(33) => 
                           state_main_out_plane0_33_port, INPUT(32) => 
                           state_main_out_plane0_32_port, INPUT(31) => 
                           state_main_out_plane0_31_port, INPUT(30) => 
                           state_main_out_plane0_30_port, INPUT(29) => 
                           state_main_out_plane0_29_port, INPUT(28) => 
                           state_main_out_plane0_28_port, INPUT(27) => 
                           state_main_out_plane0_27_port, INPUT(26) => 
                           state_main_out_plane0_26_port, INPUT(25) => 
                           state_main_out_plane0_25_port, INPUT(24) => 
                           state_main_out_plane0_24_port, INPUT(23) => 
                           state_main_out_plane0_23_port, INPUT(22) => 
                           state_main_out_plane0_22_port, INPUT(21) => 
                           state_main_out_plane0_21_port, INPUT(20) => 
                           state_main_out_plane0_20_port, INPUT(19) => 
                           state_main_out_plane0_19_port, INPUT(18) => 
                           state_main_out_plane0_18_port, INPUT(17) => 
                           state_main_out_plane0_17_port, INPUT(16) => 
                           state_main_out_plane0_16_port, INPUT(15) => 
                           state_main_out_plane0_15_port, INPUT(14) => 
                           state_main_out_plane0_14_port, INPUT(13) => 
                           state_main_out_plane0_13_port, INPUT(12) => 
                           state_main_out_plane0_12_port, INPUT(11) => 
                           state_main_out_plane0_11_port, INPUT(10) => 
                           state_main_out_plane0_10_port, INPUT(9) => 
                           state_main_out_plane0_9_port, INPUT(8) => 
                           state_main_out_plane0_8_port, INPUT(7) => 
                           state_main_out_plane0_7_port, INPUT(6) => 
                           state_main_out_plane0_6_port, INPUT(5) => 
                           state_main_out_plane0_5_port, INPUT(4) => 
                           state_main_out_plane0_4_port, INPUT(3) => 
                           state_main_out_plane0_3_port, INPUT(2) => 
                           state_main_out_plane0_2_port, INPUT(1) => 
                           state_main_out_plane0_1_port, INPUT(0) => 
                           state_main_out_plane0_0_port, perm_output(383) => 
                           perm_output_383_port, perm_output(382) => 
                           perm_output_382_port, perm_output(381) => 
                           perm_output_381_port, perm_output(380) => 
                           perm_output_380_port, perm_output(379) => 
                           perm_output_379_port, perm_output(378) => 
                           perm_output_378_port, perm_output(377) => 
                           perm_output_377_port, perm_output(376) => 
                           perm_output_376_port, perm_output(375) => 
                           perm_output_375_port, perm_output(374) => 
                           perm_output_374_port, perm_output(373) => 
                           perm_output_373_port, perm_output(372) => 
                           perm_output_372_port, perm_output(371) => 
                           perm_output_371_port, perm_output(370) => 
                           perm_output_370_port, perm_output(369) => 
                           perm_output_369_port, perm_output(368) => 
                           perm_output_368_port, perm_output(367) => 
                           perm_output_367_port, perm_output(366) => 
                           perm_output_366_port, perm_output(365) => 
                           perm_output_365_port, perm_output(364) => 
                           perm_output_364_port, perm_output(363) => 
                           perm_output_363_port, perm_output(362) => 
                           perm_output_362_port, perm_output(361) => 
                           perm_output_361_port, perm_output(360) => 
                           perm_output_360_port, perm_output(359) => 
                           perm_output_359_port, perm_output(358) => 
                           perm_output_358_port, perm_output(357) => 
                           perm_output_357_port, perm_output(356) => 
                           perm_output_356_port, perm_output(355) => 
                           perm_output_355_port, perm_output(354) => 
                           perm_output_354_port, perm_output(353) => 
                           perm_output_353_port, perm_output(352) => 
                           perm_output_352_port, perm_output(351) => 
                           perm_output_351_port, perm_output(350) => 
                           perm_output_350_port, perm_output(349) => 
                           perm_output_349_port, perm_output(348) => 
                           perm_output_348_port, perm_output(347) => 
                           perm_output_347_port, perm_output(346) => 
                           perm_output_346_port, perm_output(345) => 
                           perm_output_345_port, perm_output(344) => 
                           perm_output_344_port, perm_output(343) => 
                           perm_output_343_port, perm_output(342) => 
                           perm_output_342_port, perm_output(341) => 
                           perm_output_341_port, perm_output(340) => 
                           perm_output_340_port, perm_output(339) => 
                           perm_output_339_port, perm_output(338) => 
                           perm_output_338_port, perm_output(337) => 
                           perm_output_337_port, perm_output(336) => 
                           perm_output_336_port, perm_output(335) => 
                           perm_output_335_port, perm_output(334) => 
                           perm_output_334_port, perm_output(333) => 
                           perm_output_333_port, perm_output(332) => 
                           perm_output_332_port, perm_output(331) => 
                           perm_output_331_port, perm_output(330) => 
                           perm_output_330_port, perm_output(329) => 
                           perm_output_329_port, perm_output(328) => 
                           perm_output_328_port, perm_output(327) => 
                           perm_output_327_port, perm_output(326) => 
                           perm_output_326_port, perm_output(325) => 
                           perm_output_325_port, perm_output(324) => 
                           perm_output_324_port, perm_output(323) => 
                           perm_output_323_port, perm_output(322) => 
                           perm_output_322_port, perm_output(321) => 
                           perm_output_321_port, perm_output(320) => 
                           perm_output_320_port, perm_output(319) => 
                           perm_output_319_port, perm_output(318) => 
                           perm_output_318_port, perm_output(317) => 
                           perm_output_317_port, perm_output(316) => 
                           perm_output_316_port, perm_output(315) => 
                           perm_output_315_port, perm_output(314) => 
                           perm_output_314_port, perm_output(313) => 
                           perm_output_313_port, perm_output(312) => 
                           perm_output_312_port, perm_output(311) => 
                           perm_output_311_port, perm_output(310) => 
                           perm_output_310_port, perm_output(309) => 
                           perm_output_309_port, perm_output(308) => 
                           perm_output_308_port, perm_output(307) => 
                           perm_output_307_port, perm_output(306) => 
                           perm_output_306_port, perm_output(305) => 
                           perm_output_305_port, perm_output(304) => 
                           perm_output_304_port, perm_output(303) => 
                           perm_output_303_port, perm_output(302) => 
                           perm_output_302_port, perm_output(301) => 
                           perm_output_301_port, perm_output(300) => 
                           perm_output_300_port, perm_output(299) => 
                           perm_output_299_port, perm_output(298) => 
                           perm_output_298_port, perm_output(297) => 
                           perm_output_297_port, perm_output(296) => 
                           perm_output_296_port, perm_output(295) => 
                           perm_output_295_port, perm_output(294) => 
                           perm_output_294_port, perm_output(293) => 
                           perm_output_293_port, perm_output(292) => 
                           perm_output_292_port, perm_output(291) => 
                           perm_output_291_port, perm_output(290) => 
                           perm_output_290_port, perm_output(289) => 
                           perm_output_289_port, perm_output(288) => 
                           perm_output_288_port, perm_output(287) => 
                           perm_output_287_port, perm_output(286) => 
                           perm_output_286_port, perm_output(285) => 
                           perm_output_285_port, perm_output(284) => 
                           perm_output_284_port, perm_output(283) => 
                           perm_output_283_port, perm_output(282) => 
                           perm_output_282_port, perm_output(281) => 
                           perm_output_281_port, perm_output(280) => 
                           perm_output_280_port, perm_output(279) => 
                           perm_output_279_port, perm_output(278) => 
                           perm_output_278_port, perm_output(277) => 
                           perm_output_277_port, perm_output(276) => 
                           perm_output_276_port, perm_output(275) => 
                           perm_output_275_port, perm_output(274) => 
                           perm_output_274_port, perm_output(273) => 
                           perm_output_273_port, perm_output(272) => 
                           perm_output_272_port, perm_output(271) => 
                           perm_output_271_port, perm_output(270) => 
                           perm_output_270_port, perm_output(269) => 
                           perm_output_269_port, perm_output(268) => 
                           perm_output_268_port, perm_output(267) => 
                           perm_output_267_port, perm_output(266) => 
                           perm_output_266_port, perm_output(265) => 
                           perm_output_265_port, perm_output(264) => 
                           perm_output_264_port, perm_output(263) => 
                           perm_output_263_port, perm_output(262) => 
                           perm_output_262_port, perm_output(261) => 
                           perm_output_261_port, perm_output(260) => 
                           perm_output_260_port, perm_output(259) => 
                           perm_output_259_port, perm_output(258) => 
                           perm_output_258_port, perm_output(257) => 
                           perm_output_257_port, perm_output(256) => 
                           perm_output_256_port, perm_output(255) => 
                           perm_output_255_port, perm_output(254) => 
                           perm_output_254_port, perm_output(253) => 
                           perm_output_253_port, perm_output(252) => 
                           perm_output_252_port, perm_output(251) => 
                           perm_output_251_port, perm_output(250) => 
                           perm_output_250_port, perm_output(249) => 
                           perm_output_249_port, perm_output(248) => 
                           perm_output_248_port, perm_output(247) => 
                           perm_output_247_port, perm_output(246) => 
                           perm_output_246_port, perm_output(245) => 
                           perm_output_245_port, perm_output(244) => 
                           perm_output_244_port, perm_output(243) => 
                           perm_output_243_port, perm_output(242) => 
                           perm_output_242_port, perm_output(241) => 
                           perm_output_241_port, perm_output(240) => 
                           perm_output_240_port, perm_output(239) => 
                           perm_output_239_port, perm_output(238) => 
                           perm_output_238_port, perm_output(237) => 
                           perm_output_237_port, perm_output(236) => 
                           perm_output_236_port, perm_output(235) => 
                           perm_output_235_port, perm_output(234) => 
                           perm_output_234_port, perm_output(233) => 
                           perm_output_233_port, perm_output(232) => 
                           perm_output_232_port, perm_output(231) => 
                           perm_output_231_port, perm_output(230) => 
                           perm_output_230_port, perm_output(229) => 
                           perm_output_229_port, perm_output(228) => 
                           perm_output_228_port, perm_output(227) => 
                           perm_output_227_port, perm_output(226) => 
                           perm_output_226_port, perm_output(225) => 
                           perm_output_225_port, perm_output(224) => 
                           perm_output_224_port, perm_output(223) => 
                           perm_output_223_port, perm_output(222) => 
                           perm_output_222_port, perm_output(221) => 
                           perm_output_221_port, perm_output(220) => 
                           perm_output_220_port, perm_output(219) => 
                           perm_output_219_port, perm_output(218) => 
                           perm_output_218_port, perm_output(217) => 
                           perm_output_217_port, perm_output(216) => 
                           perm_output_216_port, perm_output(215) => 
                           perm_output_215_port, perm_output(214) => 
                           perm_output_214_port, perm_output(213) => 
                           perm_output_213_port, perm_output(212) => 
                           perm_output_212_port, perm_output(211) => 
                           perm_output_211_port, perm_output(210) => 
                           perm_output_210_port, perm_output(209) => 
                           perm_output_209_port, perm_output(208) => 
                           perm_output_208_port, perm_output(207) => 
                           perm_output_207_port, perm_output(206) => 
                           perm_output_206_port, perm_output(205) => 
                           perm_output_205_port, perm_output(204) => 
                           perm_output_204_port, perm_output(203) => 
                           perm_output_203_port, perm_output(202) => 
                           perm_output_202_port, perm_output(201) => 
                           perm_output_201_port, perm_output(200) => 
                           perm_output_200_port, perm_output(199) => 
                           perm_output_199_port, perm_output(198) => 
                           perm_output_198_port, perm_output(197) => 
                           perm_output_197_port, perm_output(196) => 
                           perm_output_196_port, perm_output(195) => 
                           perm_output_195_port, perm_output(194) => 
                           perm_output_194_port, perm_output(193) => 
                           perm_output_193_port, perm_output(192) => 
                           perm_output_192_port, perm_output(191) => 
                           perm_output_191_port, perm_output(190) => 
                           perm_output_190_port, perm_output(189) => 
                           perm_output_189_port, perm_output(188) => 
                           perm_output_188_port, perm_output(187) => 
                           perm_output_187_port, perm_output(186) => 
                           perm_output_186_port, perm_output(185) => 
                           perm_output_185_port, perm_output(184) => 
                           perm_output_184_port, perm_output(183) => 
                           perm_output_183_port, perm_output(182) => 
                           perm_output_182_port, perm_output(181) => 
                           perm_output_181_port, perm_output(180) => 
                           perm_output_180_port, perm_output(179) => 
                           perm_output_179_port, perm_output(178) => 
                           perm_output_178_port, perm_output(177) => 
                           perm_output_177_port, perm_output(176) => 
                           perm_output_176_port, perm_output(175) => 
                           perm_output_175_port, perm_output(174) => 
                           perm_output_174_port, perm_output(173) => 
                           perm_output_173_port, perm_output(172) => 
                           perm_output_172_port, perm_output(171) => 
                           perm_output_171_port, perm_output(170) => 
                           perm_output_170_port, perm_output(169) => 
                           perm_output_169_port, perm_output(168) => 
                           perm_output_168_port, perm_output(167) => 
                           perm_output_167_port, perm_output(166) => 
                           perm_output_166_port, perm_output(165) => 
                           perm_output_165_port, perm_output(164) => 
                           perm_output_164_port, perm_output(163) => 
                           perm_output_163_port, perm_output(162) => 
                           perm_output_162_port, perm_output(161) => 
                           perm_output_161_port, perm_output(160) => 
                           perm_output_160_port, perm_output(159) => 
                           perm_output_159_port, perm_output(158) => 
                           perm_output_158_port, perm_output(157) => 
                           perm_output_157_port, perm_output(156) => 
                           perm_output_156_port, perm_output(155) => 
                           perm_output_155_port, perm_output(154) => 
                           perm_output_154_port, perm_output(153) => 
                           perm_output_153_port, perm_output(152) => 
                           perm_output_152_port, perm_output(151) => 
                           perm_output_151_port, perm_output(150) => 
                           perm_output_150_port, perm_output(149) => 
                           perm_output_149_port, perm_output(148) => 
                           perm_output_148_port, perm_output(147) => 
                           perm_output_147_port, perm_output(146) => 
                           perm_output_146_port, perm_output(145) => 
                           perm_output_145_port, perm_output(144) => 
                           perm_output_144_port, perm_output(143) => 
                           perm_output_143_port, perm_output(142) => 
                           perm_output_142_port, perm_output(141) => 
                           perm_output_141_port, perm_output(140) => 
                           perm_output_140_port, perm_output(139) => 
                           perm_output_139_port, perm_output(138) => 
                           perm_output_138_port, perm_output(137) => 
                           perm_output_137_port, perm_output(136) => 
                           perm_output_136_port, perm_output(135) => 
                           perm_output_135_port, perm_output(134) => 
                           perm_output_134_port, perm_output(133) => 
                           perm_output_133_port, perm_output(132) => 
                           perm_output_132_port, perm_output(131) => 
                           perm_output_131_port, perm_output(130) => 
                           perm_output_130_port, perm_output(129) => 
                           perm_output_129_port, perm_output(128) => 
                           perm_output_128_port, perm_output(127) => 
                           perm_output_127_port, perm_output(126) => 
                           perm_output_126_port, perm_output(125) => 
                           perm_output_125_port, perm_output(124) => 
                           perm_output_124_port, perm_output(123) => 
                           perm_output_123_port, perm_output(122) => 
                           perm_output_122_port, perm_output(121) => 
                           perm_output_121_port, perm_output(120) => 
                           perm_output_120_port, perm_output(119) => 
                           perm_output_119_port, perm_output(118) => 
                           perm_output_118_port, perm_output(117) => 
                           perm_output_117_port, perm_output(116) => 
                           perm_output_116_port, perm_output(115) => 
                           perm_output_115_port, perm_output(114) => 
                           perm_output_114_port, perm_output(113) => 
                           perm_output_113_port, perm_output(112) => 
                           perm_output_112_port, perm_output(111) => 
                           perm_output_111_port, perm_output(110) => 
                           perm_output_110_port, perm_output(109) => 
                           perm_output_109_port, perm_output(108) => 
                           perm_output_108_port, perm_output(107) => 
                           perm_output_107_port, perm_output(106) => 
                           perm_output_106_port, perm_output(105) => 
                           perm_output_105_port, perm_output(104) => 
                           perm_output_104_port, perm_output(103) => 
                           perm_output_103_port, perm_output(102) => 
                           perm_output_102_port, perm_output(101) => 
                           perm_output_101_port, perm_output(100) => 
                           perm_output_100_port, perm_output(99) => 
                           perm_output_99_port, perm_output(98) => 
                           perm_output_98_port, perm_output(97) => 
                           perm_output_97_port, perm_output(96) => 
                           perm_output_96_port, perm_output(95) => 
                           perm_output_95_port, perm_output(94) => 
                           perm_output_94_port, perm_output(93) => 
                           perm_output_93_port, perm_output(92) => 
                           perm_output_92_port, perm_output(91) => 
                           perm_output_91_port, perm_output(90) => 
                           perm_output_90_port, perm_output(89) => 
                           perm_output_89_port, perm_output(88) => 
                           perm_output_88_port, perm_output(87) => 
                           perm_output_87_port, perm_output(86) => 
                           perm_output_86_port, perm_output(85) => 
                           perm_output_85_port, perm_output(84) => 
                           perm_output_84_port, perm_output(83) => 
                           perm_output_83_port, perm_output(82) => 
                           perm_output_82_port, perm_output(81) => 
                           perm_output_81_port, perm_output(80) => 
                           perm_output_80_port, perm_output(79) => 
                           perm_output_79_port, perm_output(78) => 
                           perm_output_78_port, perm_output(77) => 
                           perm_output_77_port, perm_output(76) => 
                           perm_output_76_port, perm_output(75) => 
                           perm_output_75_port, perm_output(74) => 
                           perm_output_74_port, perm_output(73) => 
                           perm_output_73_port, perm_output(72) => 
                           perm_output_72_port, perm_output(71) => 
                           perm_output_71_port, perm_output(70) => 
                           perm_output_70_port, perm_output(69) => 
                           perm_output_69_port, perm_output(68) => 
                           perm_output_68_port, perm_output(67) => 
                           perm_output_67_port, perm_output(66) => 
                           perm_output_66_port, perm_output(65) => 
                           perm_output_65_port, perm_output(64) => 
                           perm_output_64_port, perm_output(63) => 
                           perm_output_63_port, perm_output(62) => 
                           perm_output_62_port, perm_output(61) => 
                           perm_output_61_port, perm_output(60) => 
                           perm_output_60_port, perm_output(59) => 
                           perm_output_59_port, perm_output(58) => 
                           perm_output_58_port, perm_output(57) => 
                           perm_output_57_port, perm_output(56) => 
                           perm_output_56_port, perm_output(55) => 
                           perm_output_55_port, perm_output(54) => 
                           perm_output_54_port, perm_output(53) => 
                           perm_output_53_port, perm_output(52) => 
                           perm_output_52_port, perm_output(51) => 
                           perm_output_51_port, perm_output(50) => 
                           perm_output_50_port, perm_output(49) => 
                           perm_output_49_port, perm_output(48) => 
                           perm_output_48_port, perm_output(47) => 
                           perm_output_47_port, perm_output(46) => 
                           perm_output_46_port, perm_output(45) => 
                           perm_output_45_port, perm_output(44) => 
                           perm_output_44_port, perm_output(43) => 
                           perm_output_43_port, perm_output(42) => 
                           perm_output_42_port, perm_output(41) => 
                           perm_output_41_port, perm_output(40) => 
                           perm_output_40_port, perm_output(39) => 
                           perm_output_39_port, perm_output(38) => 
                           perm_output_38_port, perm_output(37) => 
                           perm_output_37_port, perm_output(36) => 
                           perm_output_36_port, perm_output(35) => 
                           perm_output_35_port, perm_output(34) => 
                           perm_output_34_port, perm_output(33) => 
                           perm_output_33_port, perm_output(32) => 
                           perm_output_32_port, perm_output(31) => 
                           perm_output_31_port, perm_output(30) => 
                           perm_output_30_port, perm_output(29) => 
                           perm_output_29_port, perm_output(28) => 
                           perm_output_28_port, perm_output(27) => 
                           perm_output_27_port, perm_output(26) => 
                           perm_output_26_port, perm_output(25) => 
                           perm_output_25_port, perm_output(24) => 
                           perm_output_24_port, perm_output(23) => 
                           perm_output_23_port, perm_output(22) => 
                           perm_output_22_port, perm_output(21) => 
                           perm_output_21_port, perm_output(20) => 
                           perm_output_20_port, perm_output(19) => 
                           perm_output_19_port, perm_output(18) => 
                           perm_output_18_port, perm_output(17) => 
                           perm_output_17_port, perm_output(16) => 
                           perm_output_16_port, perm_output(15) => 
                           perm_output_15_port, perm_output(14) => 
                           perm_output_14_port, perm_output(13) => 
                           perm_output_13_port, perm_output(12) => 
                           perm_output_12_port, perm_output(11) => 
                           perm_output_11_port, perm_output(10) => 
                           perm_output_10_port, perm_output(9) => 
                           perm_output_9_port, perm_output(8) => 
                           perm_output_8_port, perm_output(7) => 
                           perm_output_7_port, perm_output(6) => 
                           perm_output_6_port, perm_output(5) => 
                           perm_output_5_port, perm_output(4) => 
                           perm_output_4_port, perm_output(3) => 
                           perm_output_3_port, perm_output(2) => 
                           perm_output_2_port, perm_output(1) => 
                           perm_output_1_port, perm_output(0) => 
                           perm_output_0_port, RNDCTR(3) => rnd_counter(3), 
                           RNDCTR(2) => rnd_counter(2), RNDCTR(1) => 
                           rnd_counter(1), RNDCTR(0) => rnd_counter(0));
   I_0 : GTECH_NOT port map( A => extract_sel, Z => N571);
   I_1 : GTECH_NOT port map( A => xor_sel, Z => N572);
   I_2 : GTECH_NOT port map( A => cyc_state_update_sel, Z => N573);
   I_3 : GTECH_NOT port map( A => state_main_sel(6), Z => N574);
   C1634_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 128 )
      port map(
         -- Connections to port 'DATA1'
         DATA(127) => state_main_out_plane0_127_port, DATA(126) => 
               state_main_out_plane0_126_port, DATA(125) => 
               state_main_out_plane0_125_port, DATA(124) => 
               state_main_out_plane0_124_port, DATA(123) => 
               state_main_out_plane0_123_port, DATA(122) => 
               state_main_out_plane0_122_port, DATA(121) => 
               state_main_out_plane0_121_port, DATA(120) => 
               state_main_out_plane0_120_port, DATA(119) => 
               state_main_out_plane0_119_port, DATA(118) => 
               state_main_out_plane0_118_port, DATA(117) => 
               state_main_out_plane0_117_port, DATA(116) => 
               state_main_out_plane0_116_port, DATA(115) => 
               state_main_out_plane0_115_port, DATA(114) => 
               state_main_out_plane0_114_port, DATA(113) => 
               state_main_out_plane0_113_port, DATA(112) => 
               state_main_out_plane0_112_port, DATA(111) => 
               state_main_out_plane0_111_port, DATA(110) => 
               state_main_out_plane0_110_port, DATA(109) => 
               state_main_out_plane0_109_port, DATA(108) => 
               state_main_out_plane0_108_port, DATA(107) => 
               state_main_out_plane0_107_port, DATA(106) => 
               state_main_out_plane0_106_port, DATA(105) => 
               state_main_out_plane0_105_port, DATA(104) => 
               state_main_out_plane0_104_port, DATA(103) => 
               state_main_out_plane0_103_port, DATA(102) => 
               state_main_out_plane0_102_port, DATA(101) => 
               state_main_out_plane0_101_port, DATA(100) => 
               state_main_out_plane0_100_port, DATA(99) => 
               state_main_out_plane0_99_port, DATA(98) => 
               state_main_out_plane0_98_port, DATA(97) => 
               state_main_out_plane0_97_port, DATA(96) => 
               state_main_out_plane0_96_port, DATA(95) => 
               state_main_out_plane0_95_port, DATA(94) => 
               state_main_out_plane0_94_port, DATA(93) => 
               state_main_out_plane0_93_port, DATA(92) => 
               state_main_out_plane0_92_port, DATA(91) => 
               state_main_out_plane0_91_port, DATA(90) => 
               state_main_out_plane0_90_port, DATA(89) => 
               state_main_out_plane0_89_port, DATA(88) => 
               state_main_out_plane0_88_port, DATA(87) => 
               state_main_out_plane0_87_port, DATA(86) => 
               state_main_out_plane0_86_port, DATA(85) => 
               state_main_out_plane0_85_port, DATA(84) => 
               state_main_out_plane0_84_port, DATA(83) => 
               state_main_out_plane0_83_port, DATA(82) => 
               state_main_out_plane0_82_port, DATA(81) => 
               state_main_out_plane0_81_port, DATA(80) => 
               state_main_out_plane0_80_port, DATA(79) => 
               state_main_out_plane0_79_port, DATA(78) => 
               state_main_out_plane0_78_port, DATA(77) => 
               state_main_out_plane0_77_port, DATA(76) => 
               state_main_out_plane0_76_port, DATA(75) => 
               state_main_out_plane0_75_port, DATA(74) => 
               state_main_out_plane0_74_port, DATA(73) => 
               state_main_out_plane0_73_port, DATA(72) => 
               state_main_out_plane0_72_port, DATA(71) => 
               state_main_out_plane0_71_port, DATA(70) => 
               state_main_out_plane0_70_port, DATA(69) => 
               state_main_out_plane0_69_port, DATA(68) => 
               state_main_out_plane0_68_port, DATA(67) => 
               state_main_out_plane0_67_port, DATA(66) => 
               state_main_out_plane0_66_port, DATA(65) => 
               state_main_out_plane0_65_port, DATA(64) => 
               state_main_out_plane0_64_port, DATA(63) => 
               state_main_out_plane0_63_port, DATA(62) => 
               state_main_out_plane0_62_port, DATA(61) => 
               state_main_out_plane0_61_port, DATA(60) => 
               state_main_out_plane0_60_port, DATA(59) => 
               state_main_out_plane0_59_port, DATA(58) => 
               state_main_out_plane0_58_port, DATA(57) => 
               state_main_out_plane0_57_port, DATA(56) => 
               state_main_out_plane0_56_port, DATA(55) => 
               state_main_out_plane0_55_port, DATA(54) => 
               state_main_out_plane0_54_port, DATA(53) => 
               state_main_out_plane0_53_port, DATA(52) => 
               state_main_out_plane0_52_port, DATA(51) => 
               state_main_out_plane0_51_port, DATA(50) => 
               state_main_out_plane0_50_port, DATA(49) => 
               state_main_out_plane0_49_port, DATA(48) => 
               state_main_out_plane0_48_port, DATA(47) => 
               state_main_out_plane0_47_port, DATA(46) => 
               state_main_out_plane0_46_port, DATA(45) => 
               state_main_out_plane0_45_port, DATA(44) => 
               state_main_out_plane0_44_port, DATA(43) => 
               state_main_out_plane0_43_port, DATA(42) => 
               state_main_out_plane0_42_port, DATA(41) => 
               state_main_out_plane0_41_port, DATA(40) => 
               state_main_out_plane0_40_port, DATA(39) => 
               state_main_out_plane0_39_port, DATA(38) => 
               state_main_out_plane0_38_port, DATA(37) => 
               state_main_out_plane0_37_port, DATA(36) => 
               state_main_out_plane0_36_port, DATA(35) => 
               state_main_out_plane0_35_port, DATA(34) => 
               state_main_out_plane0_34_port, DATA(33) => 
               state_main_out_plane0_33_port, DATA(32) => 
               state_main_out_plane0_32_port, DATA(31) => 
               state_main_out_plane0_31_port, DATA(30) => 
               state_main_out_plane0_30_port, DATA(29) => 
               state_main_out_plane0_29_port, DATA(28) => 
               state_main_out_plane0_28_port, DATA(27) => 
               state_main_out_plane0_27_port, DATA(26) => 
               state_main_out_plane0_26_port, DATA(25) => 
               state_main_out_plane0_25_port, DATA(24) => 
               state_main_out_plane0_24_port, DATA(23) => 
               state_main_out_plane0_23_port, DATA(22) => 
               state_main_out_plane0_22_port, DATA(21) => 
               state_main_out_plane0_21_port, DATA(20) => 
               state_main_out_plane0_20_port, DATA(19) => 
               state_main_out_plane0_19_port, DATA(18) => 
               state_main_out_plane0_18_port, DATA(17) => 
               state_main_out_plane0_17_port, DATA(16) => 
               state_main_out_plane0_16_port, DATA(15) => 
               state_main_out_plane0_15_port, DATA(14) => 
               state_main_out_plane0_14_port, DATA(13) => 
               state_main_out_plane0_13_port, DATA(12) => 
               state_main_out_plane0_12_port, DATA(11) => 
               state_main_out_plane0_11_port, DATA(10) => 
               state_main_out_plane0_10_port, DATA(9) => 
               state_main_out_plane0_9_port, DATA(8) => 
               state_main_out_plane0_8_port, DATA(7) => 
               state_main_out_plane0_7_port, DATA(6) => 
               state_main_out_plane0_6_port, DATA(5) => 
               state_main_out_plane0_5_port, DATA(4) => 
               state_main_out_plane0_4_port, DATA(3) => 
               state_main_out_plane0_3_port, DATA(2) => 
               state_main_out_plane0_2_port, DATA(1) => 
               state_main_out_plane0_1_port, DATA(0) => 
               state_main_out_plane0_0_port, 
         -- Connections to port 'DATA2'
         DATA(255) => state_main_out_plane1_127_port, DATA(254) => 
               state_main_out_plane1_126_port, DATA(253) => 
               state_main_out_plane1_125_port, DATA(252) => 
               state_main_out_plane1_124_port, DATA(251) => 
               state_main_out_plane1_123_port, DATA(250) => 
               state_main_out_plane1_122_port, DATA(249) => 
               state_main_out_plane1_121_port, DATA(248) => 
               state_main_out_plane1_120_port, DATA(247) => 
               state_main_out_plane1_119_port, DATA(246) => 
               state_main_out_plane1_118_port, DATA(245) => 
               state_main_out_plane1_117_port, DATA(244) => 
               state_main_out_plane1_116_port, DATA(243) => 
               state_main_out_plane1_115_port, DATA(242) => 
               state_main_out_plane1_114_port, DATA(241) => 
               state_main_out_plane1_113_port, DATA(240) => 
               state_main_out_plane1_112_port, DATA(239) => 
               state_main_out_plane1_111_port, DATA(238) => 
               state_main_out_plane1_110_port, DATA(237) => 
               state_main_out_plane1_109_port, DATA(236) => 
               state_main_out_plane1_108_port, DATA(235) => 
               state_main_out_plane1_107_port, DATA(234) => 
               state_main_out_plane1_106_port, DATA(233) => 
               state_main_out_plane1_105_port, DATA(232) => 
               state_main_out_plane1_104_port, DATA(231) => 
               state_main_out_plane1_103_port, DATA(230) => 
               state_main_out_plane1_102_port, DATA(229) => 
               state_main_out_plane1_101_port, DATA(228) => 
               state_main_out_plane1_100_port, DATA(227) => 
               state_main_out_plane1_99_port, DATA(226) => 
               state_main_out_plane1_98_port, DATA(225) => 
               state_main_out_plane1_97_port, DATA(224) => 
               state_main_out_plane1_96_port, DATA(223) => 
               state_main_out_plane1_95_port, DATA(222) => 
               state_main_out_plane1_94_port, DATA(221) => 
               state_main_out_plane1_93_port, DATA(220) => 
               state_main_out_plane1_92_port, DATA(219) => 
               state_main_out_plane1_91_port, DATA(218) => 
               state_main_out_plane1_90_port, DATA(217) => 
               state_main_out_plane1_89_port, DATA(216) => 
               state_main_out_plane1_88_port, DATA(215) => 
               state_main_out_plane1_87_port, DATA(214) => 
               state_main_out_plane1_86_port, DATA(213) => 
               state_main_out_plane1_85_port, DATA(212) => 
               state_main_out_plane1_84_port, DATA(211) => 
               state_main_out_plane1_83_port, DATA(210) => 
               state_main_out_plane1_82_port, DATA(209) => 
               state_main_out_plane1_81_port, DATA(208) => 
               state_main_out_plane1_80_port, DATA(207) => 
               state_main_out_plane1_79_port, DATA(206) => 
               state_main_out_plane1_78_port, DATA(205) => 
               state_main_out_plane1_77_port, DATA(204) => 
               state_main_out_plane1_76_port, DATA(203) => 
               state_main_out_plane1_75_port, DATA(202) => 
               state_main_out_plane1_74_port, DATA(201) => 
               state_main_out_plane1_73_port, DATA(200) => 
               state_main_out_plane1_72_port, DATA(199) => 
               state_main_out_plane1_71_port, DATA(198) => 
               state_main_out_plane1_70_port, DATA(197) => 
               state_main_out_plane1_69_port, DATA(196) => 
               state_main_out_plane1_68_port, DATA(195) => 
               state_main_out_plane1_67_port, DATA(194) => 
               state_main_out_plane1_66_port, DATA(193) => 
               state_main_out_plane1_65_port, DATA(192) => 
               state_main_out_plane1_64_port, DATA(191) => 
               state_main_out_plane1_63_port, DATA(190) => 
               state_main_out_plane1_62_port, DATA(189) => 
               state_main_out_plane1_61_port, DATA(188) => 
               state_main_out_plane1_60_port, DATA(187) => 
               state_main_out_plane1_59_port, DATA(186) => 
               state_main_out_plane1_58_port, DATA(185) => 
               state_main_out_plane1_57_port, DATA(184) => 
               state_main_out_plane1_56_port, DATA(183) => 
               state_main_out_plane1_55_port, DATA(182) => 
               state_main_out_plane1_54_port, DATA(181) => 
               state_main_out_plane1_53_port, DATA(180) => 
               state_main_out_plane1_52_port, DATA(179) => 
               state_main_out_plane1_51_port, DATA(178) => 
               state_main_out_plane1_50_port, DATA(177) => 
               state_main_out_plane1_49_port, DATA(176) => 
               state_main_out_plane1_48_port, DATA(175) => 
               state_main_out_plane1_47_port, DATA(174) => 
               state_main_out_plane1_46_port, DATA(173) => 
               state_main_out_plane1_45_port, DATA(172) => 
               state_main_out_plane1_44_port, DATA(171) => 
               state_main_out_plane1_43_port, DATA(170) => 
               state_main_out_plane1_42_port, DATA(169) => 
               state_main_out_plane1_41_port, DATA(168) => 
               state_main_out_plane1_40_port, DATA(167) => 
               state_main_out_plane1_39_port, DATA(166) => 
               state_main_out_plane1_38_port, DATA(165) => 
               state_main_out_plane1_37_port, DATA(164) => 
               state_main_out_plane1_36_port, DATA(163) => 
               state_main_out_plane1_35_port, DATA(162) => 
               state_main_out_plane1_34_port, DATA(161) => 
               state_main_out_plane1_33_port, DATA(160) => 
               state_main_out_plane1_32_port, DATA(159) => 
               state_main_out_plane1_31_port, DATA(158) => 
               state_main_out_plane1_30_port, DATA(157) => 
               state_main_out_plane1_29_port, DATA(156) => 
               state_main_out_plane1_28_port, DATA(155) => 
               state_main_out_plane1_27_port, DATA(154) => 
               state_main_out_plane1_26_port, DATA(153) => 
               state_main_out_plane1_25_port, DATA(152) => 
               state_main_out_plane1_24_port, DATA(151) => 
               state_main_out_plane1_23_port, DATA(150) => 
               state_main_out_plane1_22_port, DATA(149) => 
               state_main_out_plane1_21_port, DATA(148) => 
               state_main_out_plane1_20_port, DATA(147) => 
               state_main_out_plane1_19_port, DATA(146) => 
               state_main_out_plane1_18_port, DATA(145) => 
               state_main_out_plane1_17_port, DATA(144) => 
               state_main_out_plane1_16_port, DATA(143) => 
               state_main_out_plane1_15_port, DATA(142) => 
               state_main_out_plane1_14_port, DATA(141) => 
               state_main_out_plane1_13_port, DATA(140) => 
               state_main_out_plane1_12_port, DATA(139) => 
               state_main_out_plane1_11_port, DATA(138) => 
               state_main_out_plane1_10_port, DATA(137) => 
               state_main_out_plane1_9_port, DATA(136) => 
               state_main_out_plane1_8_port, DATA(135) => 
               state_main_out_plane1_7_port, DATA(134) => 
               state_main_out_plane1_6_port, DATA(133) => 
               state_main_out_plane1_5_port, DATA(132) => 
               state_main_out_plane1_4_port, DATA(131) => 
               state_main_out_plane1_3_port, DATA(130) => 
               state_main_out_plane1_2_port, DATA(129) => 
               state_main_out_plane1_1_port, DATA(128) => 
               state_main_out_plane1_0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N0, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N1, 
         -- Connections to port 'Z'
         Z(127) => N161, Z(126) => N160, Z(125) => N159, Z(124) => N158, Z(123)
               => N157, Z(122) => N156, Z(121) => N155, Z(120) => N154, Z(119) 
               => N153, Z(118) => N152, Z(117) => N151, Z(116) => N150, Z(115) 
               => N149, Z(114) => N148, Z(113) => N147, Z(112) => N146, Z(111) 
               => N145, Z(110) => N144, Z(109) => N143, Z(108) => N142, Z(107) 
               => N141, Z(106) => N140, Z(105) => N139, Z(104) => N138, Z(103) 
               => N137, Z(102) => N136, Z(101) => N135, Z(100) => N134, Z(99) 
               => N133, Z(98) => N132, Z(97) => N131, Z(96) => N130, Z(95) => 
               N129, Z(94) => N128, Z(93) => N127, Z(92) => N126, Z(91) => N125
               , Z(90) => N124, Z(89) => N123, Z(88) => N122, Z(87) => N121, 
               Z(86) => N120, Z(85) => N119, Z(84) => N118, Z(83) => N117, 
               Z(82) => N116, Z(81) => N115, Z(80) => N114, Z(79) => N113, 
               Z(78) => N112, Z(77) => N111, Z(76) => N110, Z(75) => N109, 
               Z(74) => N108, Z(73) => N107, Z(72) => N106, Z(71) => N105, 
               Z(70) => N104, Z(69) => N103, Z(68) => N102, Z(67) => N101, 
               Z(66) => N100, Z(65) => N99, Z(64) => N98, Z(63) => N97, Z(62) 
               => N96, Z(61) => N95, Z(60) => N94, Z(59) => N93, Z(58) => N92, 
               Z(57) => N91, Z(56) => N90, Z(55) => N89, Z(54) => N88, Z(53) =>
               N87, Z(52) => N86, Z(51) => N85, Z(50) => N84, Z(49) => N83, 
               Z(48) => N82, Z(47) => N81, Z(46) => N80, Z(45) => N79, Z(44) =>
               N78, Z(43) => N77, Z(42) => N76, Z(41) => N75, Z(40) => N74, 
               Z(39) => N73, Z(38) => N72, Z(37) => N71, Z(36) => N70, Z(35) =>
               N69, Z(34) => N68, Z(33) => N67, Z(32) => N66, Z(31) => N65, 
               Z(30) => N64, Z(29) => N63, Z(28) => N62, Z(27) => N61, Z(26) =>
               N60, Z(25) => N59, Z(24) => N58, Z(23) => N57, Z(22) => N56, 
               Z(21) => N55, Z(20) => N54, Z(19) => N53, Z(18) => N52, Z(17) =>
               N51, Z(16) => N50, Z(15) => N49, Z(14) => N48, Z(13) => N47, 
               Z(12) => N46, Z(11) => N45, Z(10) => N44, Z(9) => N43, Z(8) => 
               N42, Z(7) => N41, Z(6) => N40, Z(5) => N39, Z(4) => N38, Z(3) =>
               N37, Z(2) => N36, Z(1) => N35, Z(0) => N34 );
   B_0 : GTECH_BUF port map( A => N33, Z => N0);
   B_1 : GTECH_BUF port map( A => dcount_in(2), Z => N1);
   C1635_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 128 )
      port map(
         -- Connections to port 'DATA1'
         DATA(127) => N161, DATA(126) => N160, DATA(125) => N159, DATA(124) => 
               N158, DATA(123) => N157, DATA(122) => N156, DATA(121) => N155, 
               DATA(120) => N154, DATA(119) => N153, DATA(118) => N152, 
               DATA(117) => N151, DATA(116) => N150, DATA(115) => N149, 
               DATA(114) => N148, DATA(113) => N147, DATA(112) => N146, 
               DATA(111) => N145, DATA(110) => N144, DATA(109) => N143, 
               DATA(108) => N142, DATA(107) => N141, DATA(106) => N140, 
               DATA(105) => N139, DATA(104) => N138, DATA(103) => N137, 
               DATA(102) => N136, DATA(101) => N135, DATA(100) => N134, 
               DATA(99) => N133, DATA(98) => N132, DATA(97) => N131, DATA(96) 
               => N130, DATA(95) => N129, DATA(94) => N128, DATA(93) => N127, 
               DATA(92) => N126, DATA(91) => N125, DATA(90) => N124, DATA(89) 
               => N123, DATA(88) => N122, DATA(87) => N121, DATA(86) => N120, 
               DATA(85) => N119, DATA(84) => N118, DATA(83) => N117, DATA(82) 
               => N116, DATA(81) => N115, DATA(80) => N114, DATA(79) => N113, 
               DATA(78) => N112, DATA(77) => N111, DATA(76) => N110, DATA(75) 
               => N109, DATA(74) => N108, DATA(73) => N107, DATA(72) => N106, 
               DATA(71) => N105, DATA(70) => N104, DATA(69) => N103, DATA(68) 
               => N102, DATA(67) => N101, DATA(66) => N100, DATA(65) => N99, 
               DATA(64) => N98, DATA(63) => N97, DATA(62) => N96, DATA(61) => 
               N95, DATA(60) => N94, DATA(59) => N93, DATA(58) => N92, DATA(57)
               => N91, DATA(56) => N90, DATA(55) => N89, DATA(54) => N88, 
               DATA(53) => N87, DATA(52) => N86, DATA(51) => N85, DATA(50) => 
               N84, DATA(49) => N83, DATA(48) => N82, DATA(47) => N81, DATA(46)
               => N80, DATA(45) => N79, DATA(44) => N78, DATA(43) => N77, 
               DATA(42) => N76, DATA(41) => N75, DATA(40) => N74, DATA(39) => 
               N73, DATA(38) => N72, DATA(37) => N71, DATA(36) => N70, DATA(35)
               => N69, DATA(34) => N68, DATA(33) => N67, DATA(32) => N66, 
               DATA(31) => N65, DATA(30) => N64, DATA(29) => N63, DATA(28) => 
               N62, DATA(27) => N61, DATA(26) => N60, DATA(25) => N59, DATA(24)
               => N58, DATA(23) => N57, DATA(22) => N56, DATA(21) => N55, 
               DATA(20) => N54, DATA(19) => N53, DATA(18) => N52, DATA(17) => 
               N51, DATA(16) => N50, DATA(15) => N49, DATA(14) => N48, DATA(13)
               => N47, DATA(12) => N46, DATA(11) => N45, DATA(10) => N44, 
               DATA(9) => N43, DATA(8) => N42, DATA(7) => N41, DATA(6) => N40, 
               DATA(5) => N39, DATA(4) => N38, DATA(3) => N37, DATA(2) => N36, 
               DATA(1) => N35, DATA(0) => N34, 
         -- Connections to port 'DATA2'
         DATA(255) => state_main_out_plane2_127_port, DATA(254) => 
               state_main_out_plane2_126_port, DATA(253) => 
               state_main_out_plane2_125_port, DATA(252) => 
               state_main_out_plane2_124_port, DATA(251) => 
               state_main_out_plane2_123_port, DATA(250) => 
               state_main_out_plane2_122_port, DATA(249) => 
               state_main_out_plane2_121_port, DATA(248) => 
               state_main_out_plane2_120_port, DATA(247) => 
               state_main_out_plane2_119_port, DATA(246) => 
               state_main_out_plane2_118_port, DATA(245) => 
               state_main_out_plane2_117_port, DATA(244) => 
               state_main_out_plane2_116_port, DATA(243) => 
               state_main_out_plane2_115_port, DATA(242) => 
               state_main_out_plane2_114_port, DATA(241) => 
               state_main_out_plane2_113_port, DATA(240) => 
               state_main_out_plane2_112_port, DATA(239) => 
               state_main_out_plane2_111_port, DATA(238) => 
               state_main_out_plane2_110_port, DATA(237) => 
               state_main_out_plane2_109_port, DATA(236) => 
               state_main_out_plane2_108_port, DATA(235) => 
               state_main_out_plane2_107_port, DATA(234) => 
               state_main_out_plane2_106_port, DATA(233) => 
               state_main_out_plane2_105_port, DATA(232) => 
               state_main_out_plane2_104_port, DATA(231) => 
               state_main_out_plane2_103_port, DATA(230) => 
               state_main_out_plane2_102_port, DATA(229) => 
               state_main_out_plane2_101_port, DATA(228) => 
               state_main_out_plane2_100_port, DATA(227) => 
               state_main_out_plane2_99_port, DATA(226) => 
               state_main_out_plane2_98_port, DATA(225) => 
               state_main_out_plane2_97_port, DATA(224) => 
               state_main_out_plane2_96_port, DATA(223) => 
               state_main_out_plane2_95_port, DATA(222) => 
               state_main_out_plane2_94_port, DATA(221) => 
               state_main_out_plane2_93_port, DATA(220) => 
               state_main_out_plane2_92_port, DATA(219) => 
               state_main_out_plane2_91_port, DATA(218) => 
               state_main_out_plane2_90_port, DATA(217) => 
               state_main_out_plane2_89_port, DATA(216) => 
               state_main_out_plane2_88_port, DATA(215) => 
               state_main_out_plane2_87_port, DATA(214) => 
               state_main_out_plane2_86_port, DATA(213) => 
               state_main_out_plane2_85_port, DATA(212) => 
               state_main_out_plane2_84_port, DATA(211) => 
               state_main_out_plane2_83_port, DATA(210) => 
               state_main_out_plane2_82_port, DATA(209) => 
               state_main_out_plane2_81_port, DATA(208) => 
               state_main_out_plane2_80_port, DATA(207) => 
               state_main_out_plane2_79_port, DATA(206) => 
               state_main_out_plane2_78_port, DATA(205) => 
               state_main_out_plane2_77_port, DATA(204) => 
               state_main_out_plane2_76_port, DATA(203) => 
               state_main_out_plane2_75_port, DATA(202) => 
               state_main_out_plane2_74_port, DATA(201) => 
               state_main_out_plane2_73_port, DATA(200) => 
               state_main_out_plane2_72_port, DATA(199) => 
               state_main_out_plane2_71_port, DATA(198) => 
               state_main_out_plane2_70_port, DATA(197) => 
               state_main_out_plane2_69_port, DATA(196) => 
               state_main_out_plane2_68_port, DATA(195) => 
               state_main_out_plane2_67_port, DATA(194) => 
               state_main_out_plane2_66_port, DATA(193) => 
               state_main_out_plane2_65_port, DATA(192) => 
               state_main_out_plane2_64_port, DATA(191) => 
               state_main_out_plane2_63_port, DATA(190) => 
               state_main_out_plane2_62_port, DATA(189) => 
               state_main_out_plane2_61_port, DATA(188) => 
               state_main_out_plane2_60_port, DATA(187) => 
               state_main_out_plane2_59_port, DATA(186) => 
               state_main_out_plane2_58_port, DATA(185) => 
               state_main_out_plane2_57_port, DATA(184) => 
               state_main_out_plane2_56_port, DATA(183) => 
               state_main_out_plane2_55_port, DATA(182) => 
               state_main_out_plane2_54_port, DATA(181) => 
               state_main_out_plane2_53_port, DATA(180) => 
               state_main_out_plane2_52_port, DATA(179) => 
               state_main_out_plane2_51_port, DATA(178) => 
               state_main_out_plane2_50_port, DATA(177) => 
               state_main_out_plane2_49_port, DATA(176) => 
               state_main_out_plane2_48_port, DATA(175) => 
               state_main_out_plane2_47_port, DATA(174) => 
               state_main_out_plane2_46_port, DATA(173) => 
               state_main_out_plane2_45_port, DATA(172) => 
               state_main_out_plane2_44_port, DATA(171) => 
               state_main_out_plane2_43_port, DATA(170) => 
               state_main_out_plane2_42_port, DATA(169) => 
               state_main_out_plane2_41_port, DATA(168) => 
               state_main_out_plane2_40_port, DATA(167) => 
               state_main_out_plane2_39_port, DATA(166) => 
               state_main_out_plane2_38_port, DATA(165) => 
               state_main_out_plane2_37_port, DATA(164) => 
               state_main_out_plane2_36_port, DATA(163) => 
               state_main_out_plane2_35_port, DATA(162) => 
               state_main_out_plane2_34_port, DATA(161) => 
               state_main_out_plane2_33_port, DATA(160) => 
               state_main_out_plane2_32_port, DATA(159) => 
               state_main_out_plane2_31_port, DATA(158) => 
               state_main_out_plane2_30_port, DATA(157) => 
               state_main_out_plane2_29_port, DATA(156) => 
               state_main_out_plane2_28_port, DATA(155) => 
               state_main_out_plane2_27_port, DATA(154) => 
               state_main_out_plane2_26_port, DATA(153) => 
               state_main_out_plane2_25_port, DATA(152) => 
               state_main_out_plane2_24_port, DATA(151) => 
               state_main_out_plane2_23_port, DATA(150) => 
               state_main_out_plane2_22_port, DATA(149) => 
               state_main_out_plane2_21_port, DATA(148) => 
               state_main_out_plane2_20_port, DATA(147) => 
               state_main_out_plane2_19_port, DATA(146) => 
               state_main_out_plane2_18_port, DATA(145) => 
               state_main_out_plane2_17_port, DATA(144) => 
               state_main_out_plane2_16_port, DATA(143) => 
               state_main_out_plane2_15_port, DATA(142) => 
               state_main_out_plane2_14_port, DATA(141) => 
               state_main_out_plane2_13_port, DATA(140) => 
               state_main_out_plane2_12_port, DATA(139) => 
               state_main_out_plane2_11_port, DATA(138) => 
               state_main_out_plane2_10_port, DATA(137) => 
               state_main_out_plane2_9_port, DATA(136) => 
               state_main_out_plane2_8_port, DATA(135) => 
               state_main_out_plane2_7_port, DATA(134) => 
               state_main_out_plane2_6_port, DATA(133) => 
               state_main_out_plane2_5_port, DATA(132) => 
               state_main_out_plane2_4_port, DATA(131) => 
               state_main_out_plane2_3_port, DATA(130) => 
               state_main_out_plane2_2_port, DATA(129) => 
               state_main_out_plane2_1_port, DATA(128) => 
               state_main_out_plane2_0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N2, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N3, 
         -- Connections to port 'Z'
         Z(127) => plane_x_127_port, Z(126) => plane_x_126_port, Z(125) => 
               plane_x_125_port, Z(124) => plane_x_124_port, Z(123) => 
               plane_x_123_port, Z(122) => plane_x_122_port, Z(121) => 
               plane_x_121_port, Z(120) => plane_x_120_port, Z(119) => 
               plane_x_119_port, Z(118) => plane_x_118_port, Z(117) => 
               plane_x_117_port, Z(116) => plane_x_116_port, Z(115) => 
               plane_x_115_port, Z(114) => plane_x_114_port, Z(113) => 
               plane_x_113_port, Z(112) => plane_x_112_port, Z(111) => 
               plane_x_111_port, Z(110) => plane_x_110_port, Z(109) => 
               plane_x_109_port, Z(108) => plane_x_108_port, Z(107) => 
               plane_x_107_port, Z(106) => plane_x_106_port, Z(105) => 
               plane_x_105_port, Z(104) => plane_x_104_port, Z(103) => 
               plane_x_103_port, Z(102) => plane_x_102_port, Z(101) => 
               plane_x_101_port, Z(100) => plane_x_100_port, Z(99) => 
               plane_x_99_port, Z(98) => plane_x_98_port, Z(97) => 
               plane_x_97_port, Z(96) => plane_x_96_port, Z(95) => 
               plane_x_95_port, Z(94) => plane_x_94_port, Z(93) => 
               plane_x_93_port, Z(92) => plane_x_92_port, Z(91) => 
               plane_x_91_port, Z(90) => plane_x_90_port, Z(89) => 
               plane_x_89_port, Z(88) => plane_x_88_port, Z(87) => 
               plane_x_87_port, Z(86) => plane_x_86_port, Z(85) => 
               plane_x_85_port, Z(84) => plane_x_84_port, Z(83) => 
               plane_x_83_port, Z(82) => plane_x_82_port, Z(81) => 
               plane_x_81_port, Z(80) => plane_x_80_port, Z(79) => 
               plane_x_79_port, Z(78) => plane_x_78_port, Z(77) => 
               plane_x_77_port, Z(76) => plane_x_76_port, Z(75) => 
               plane_x_75_port, Z(74) => plane_x_74_port, Z(73) => 
               plane_x_73_port, Z(72) => plane_x_72_port, Z(71) => 
               plane_x_71_port, Z(70) => plane_x_70_port, Z(69) => 
               plane_x_69_port, Z(68) => plane_x_68_port, Z(67) => 
               plane_x_67_port, Z(66) => plane_x_66_port, Z(65) => 
               plane_x_65_port, Z(64) => plane_x_64_port, Z(63) => 
               plane_x_63_port, Z(62) => plane_x_62_port, Z(61) => 
               plane_x_61_port, Z(60) => plane_x_60_port, Z(59) => 
               plane_x_59_port, Z(58) => plane_x_58_port, Z(57) => 
               plane_x_57_port, Z(56) => plane_x_56_port, Z(55) => 
               plane_x_55_port, Z(54) => plane_x_54_port, Z(53) => 
               plane_x_53_port, Z(52) => plane_x_52_port, Z(51) => 
               plane_x_51_port, Z(50) => plane_x_50_port, Z(49) => 
               plane_x_49_port, Z(48) => plane_x_48_port, Z(47) => 
               plane_x_47_port, Z(46) => plane_x_46_port, Z(45) => 
               plane_x_45_port, Z(44) => plane_x_44_port, Z(43) => 
               plane_x_43_port, Z(42) => plane_x_42_port, Z(41) => 
               plane_x_41_port, Z(40) => plane_x_40_port, Z(39) => 
               plane_x_39_port, Z(38) => plane_x_38_port, Z(37) => 
               plane_x_37_port, Z(36) => plane_x_36_port, Z(35) => 
               plane_x_35_port, Z(34) => plane_x_34_port, Z(33) => 
               plane_x_33_port, Z(32) => plane_x_32_port, Z(31) => 
               plane_x_31_port, Z(30) => plane_x_30_port, Z(29) => 
               plane_x_29_port, Z(28) => plane_x_28_port, Z(27) => 
               plane_x_27_port, Z(26) => plane_x_26_port, Z(25) => 
               plane_x_25_port, Z(24) => plane_x_24_port, Z(23) => 
               plane_x_23_port, Z(22) => plane_x_22_port, Z(21) => 
               plane_x_21_port, Z(20) => plane_x_20_port, Z(19) => 
               plane_x_19_port, Z(18) => plane_x_18_port, Z(17) => 
               plane_x_17_port, Z(16) => plane_x_16_port, Z(15) => 
               plane_x_15_port, Z(14) => plane_x_14_port, Z(13) => 
               plane_x_13_port, Z(12) => plane_x_12_port, Z(11) => 
               plane_x_11_port, Z(10) => plane_x_10_port, Z(9) => 
               plane_x_9_port, Z(8) => plane_x_8_port, Z(7) => plane_x_7_port, 
               Z(6) => plane_x_6_port, Z(5) => plane_x_5_port, Z(4) => 
               plane_x_4_port, Z(3) => plane_x_3_port, Z(2) => plane_x_2_port, 
               Z(1) => plane_x_1_port, Z(0) => plane_x_0_port );
   B_2 : GTECH_BUF port map( A => N32, Z => N2);
   B_3 : GTECH_BUF port map( A => dcount_in(3), Z => N3);
   C1636_cell : SELECT_OP
      generic map ( num_inputs => 4, input_width => 25 )
      port map(
         -- Connections to port 'DATA1'
         DATA(24) => X_Logic0_port, DATA(23) => X_Logic0_port, DATA(22) => 
               X_Logic0_port, DATA(21) => X_Logic0_port, DATA(20) => 
               X_Logic0_port, DATA(19) => X_Logic0_port, DATA(18) => 
               X_Logic0_port, DATA(17) => X_Logic0_port, DATA(16) => 
               X_Logic0_port, DATA(15) => X_Logic0_port, DATA(14) => 
               X_Logic0_port, DATA(13) => X_Logic0_port, DATA(12) => 
               X_Logic0_port, DATA(11) => X_Logic0_port, DATA(10) => 
               X_Logic0_port, DATA(9) => X_Logic0_port, DATA(8) => 
               X_Logic1_port, DATA(7) => bdi_key_31_port, DATA(6) => 
               bdi_key_30_port, DATA(5) => bdi_key_29_port, DATA(4) => 
               bdi_key_28_port, DATA(3) => bdi_key_27_port, DATA(2) => 
               bdi_key_26_port, DATA(1) => bdi_key_25_port, DATA(0) => 
               bdi_key_24_port, 
         -- Connections to port 'DATA2'
         DATA(49) => X_Logic0_port, DATA(48) => X_Logic0_port, DATA(47) => 
               X_Logic0_port, DATA(46) => X_Logic0_port, DATA(45) => 
               X_Logic0_port, DATA(44) => X_Logic0_port, DATA(43) => 
               X_Logic0_port, DATA(42) => X_Logic0_port, DATA(41) => 
               X_Logic1_port, DATA(40) => bdi_key_23_port, DATA(39) => 
               bdi_key_22_port, DATA(38) => bdi_key_21_port, DATA(37) => 
               bdi_key_20_port, DATA(36) => bdi_key_19_port, DATA(35) => 
               bdi_key_18_port, DATA(34) => bdi_key_17_port, DATA(33) => 
               bdi_key_16_port, DATA(32) => bdi_key_31_port, DATA(31) => 
               bdi_key_30_port, DATA(30) => bdi_key_29_port, DATA(29) => 
               bdi_key_28_port, DATA(28) => bdi_key_27_port, DATA(27) => 
               bdi_key_26_port, DATA(26) => bdi_key_25_port, DATA(25) => 
               bdi_key_24_port, 
         -- Connections to port 'DATA3'
         DATA(74) => X_Logic1_port, DATA(73) => bdi_key_15_port, DATA(72) => 
               bdi_key_14_port, DATA(71) => bdi_key_13_port, DATA(70) => 
               bdi_key_12_port, DATA(69) => bdi_key_11_port, DATA(68) => 
               bdi_key_10_port, DATA(67) => bdi_key_9_port, DATA(66) => 
               bdi_key_8_port, DATA(65) => bdi_key_23_port, DATA(64) => 
               bdi_key_22_port, DATA(63) => bdi_key_21_port, DATA(62) => 
               bdi_key_20_port, DATA(61) => bdi_key_19_port, DATA(60) => 
               bdi_key_18_port, DATA(59) => bdi_key_17_port, DATA(58) => 
               bdi_key_16_port, DATA(57) => bdi_key_31_port, DATA(56) => 
               bdi_key_30_port, DATA(55) => bdi_key_29_port, DATA(54) => 
               bdi_key_28_port, DATA(53) => bdi_key_27_port, DATA(52) => 
               bdi_key_26_port, DATA(51) => bdi_key_25_port, DATA(50) => 
               bdi_key_24_port, 
         -- Connections to port 'DATA4'
         DATA(99) => X_Logic0_port, DATA(98) => X_Logic0_port, DATA(97) => 
               X_Logic0_port, DATA(96) => X_Logic0_port, DATA(95) => 
               X_Logic0_port, DATA(94) => X_Logic0_port, DATA(93) => 
               X_Logic0_port, DATA(92) => X_Logic0_port, DATA(91) => 
               X_Logic0_port, DATA(90) => X_Logic0_port, DATA(89) => 
               X_Logic0_port, DATA(88) => X_Logic0_port, DATA(87) => 
               X_Logic0_port, DATA(86) => X_Logic0_port, DATA(85) => 
               X_Logic0_port, DATA(84) => X_Logic0_port, DATA(83) => 
               X_Logic0_port, DATA(82) => X_Logic0_port, DATA(81) => 
               X_Logic0_port, DATA(80) => X_Logic0_port, DATA(79) => 
               X_Logic0_port, DATA(78) => X_Logic0_port, DATA(77) => 
               X_Logic0_port, DATA(76) => X_Logic0_port, DATA(75) => 
               X_Logic1_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N4, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N5, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N6, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N7, 
         -- Connections to port 'Z'
         Z(24) => cycd_add_24_port, Z(23) => cycd_add_23_port, Z(22) => 
               cycd_add_22_port, Z(21) => cycd_add_21_port, Z(20) => 
               cycd_add_20_port, Z(19) => cycd_add_19_port, Z(18) => 
               cycd_add_18_port, Z(17) => cycd_add_17_port, Z(16) => 
               cycd_add_16_port, Z(15) => cycd_add_15_port, Z(14) => 
               cycd_add_14_port, Z(13) => cycd_add_13_port, Z(12) => 
               cycd_add_12_port, Z(11) => cycd_add_11_port, Z(10) => 
               cycd_add_10_port, Z(9) => cycd_add_9_port, Z(8) => 
               cycd_add_8_port, Z(7) => cycd_add_7_port, Z(6) => 
               cycd_add_6_port, Z(5) => cycd_add_5_port, Z(4) => 
               cycd_add_4_port, Z(3) => cycd_add_3_port, Z(2) => 
               cycd_add_2_port, Z(1) => cycd_add_1_port, Z(0) => 
               cycd_add_0_port );
   B_4 : GTECH_BUF port map( A => N163, Z => N4);
   B_5 : GTECH_BUF port map( A => N165, Z => N5);
   B_6 : GTECH_BUF port map( A => N166, Z => N6);
   B_7 : GTECH_BUF port map( A => N169, Z => N7);
   C1637_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 32 )
      port map(
         -- Connections to port 'DATA1'
         DATA(31) => bdi_key_7_port, DATA(30) => bdi_key_6_port, DATA(29) => 
               bdi_key_5_port, DATA(28) => bdi_key_4_port, DATA(27) => 
               bdi_key_3_port, DATA(26) => bdi_key_2_port, DATA(25) => 
               bdi_key_1_port, DATA(24) => bdi_key_0_port, DATA(23) => 
               bdi_key_15_port, DATA(22) => bdi_key_14_port, DATA(21) => 
               bdi_key_13_port, DATA(20) => bdi_key_12_port, DATA(19) => 
               bdi_key_11_port, DATA(18) => bdi_key_10_port, DATA(17) => 
               bdi_key_9_port, DATA(16) => bdi_key_8_port, DATA(15) => 
               bdi_key_23_port, DATA(14) => bdi_key_22_port, DATA(13) => 
               bdi_key_21_port, DATA(12) => bdi_key_20_port, DATA(11) => 
               bdi_key_19_port, DATA(10) => bdi_key_18_port, DATA(9) => 
               bdi_key_17_port, DATA(8) => bdi_key_16_port, DATA(7) => 
               bdi_key_31_port, DATA(6) => bdi_key_30_port, DATA(5) => 
               bdi_key_29_port, DATA(4) => bdi_key_28_port, DATA(3) => 
               bdi_key_27_port, DATA(2) => bdi_key_26_port, DATA(1) => 
               bdi_key_25_port, DATA(0) => bdi_key_24_port, 
         -- Connections to port 'DATA2'
         DATA(63) => X_Logic0_port, DATA(62) => X_Logic0_port, DATA(61) => 
               X_Logic0_port, DATA(60) => X_Logic0_port, DATA(59) => 
               X_Logic0_port, DATA(58) => X_Logic0_port, DATA(57) => 
               X_Logic0_port, DATA(56) => cycd_add_24_port, DATA(55) => 
               cycd_add_23_port, DATA(54) => cycd_add_22_port, DATA(53) => 
               cycd_add_21_port, DATA(52) => cycd_add_20_port, DATA(51) => 
               cycd_add_19_port, DATA(50) => cycd_add_18_port, DATA(49) => 
               cycd_add_17_port, DATA(48) => cycd_add_16_port, DATA(47) => 
               cycd_add_15_port, DATA(46) => cycd_add_14_port, DATA(45) => 
               cycd_add_13_port, DATA(44) => cycd_add_12_port, DATA(43) => 
               cycd_add_11_port, DATA(42) => cycd_add_10_port, DATA(41) => 
               cycd_add_9_port, DATA(40) => cycd_add_8_port, DATA(39) => 
               cycd_add_7_port, DATA(38) => cycd_add_6_port, DATA(37) => 
               cycd_add_5_port, DATA(36) => cycd_add_4_port, DATA(35) => 
               cycd_add_3_port, DATA(34) => cycd_add_2_port, DATA(33) => 
               cycd_add_1_port, DATA(32) => cycd_add_0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N8, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N9, 
         -- Connections to port 'Z'
         Z(31) => xor_mux_o_31_port, Z(30) => xor_mux_o_30_port, Z(29) => 
               xor_mux_o_29_port, Z(28) => xor_mux_o_28_port, Z(27) => 
               xor_mux_o_27_port, Z(26) => xor_mux_o_26_port, Z(25) => 
               xor_mux_o_25_port, Z(24) => xor_mux_o_24_port, Z(23) => 
               xor_mux_o_23_port, Z(22) => xor_mux_o_22_port, Z(21) => 
               xor_mux_o_21_port, Z(20) => xor_mux_o_20_port, Z(19) => 
               xor_mux_o_19_port, Z(18) => xor_mux_o_18_port, Z(17) => 
               xor_mux_o_17_port, Z(16) => xor_mux_o_16_port, Z(15) => 
               xor_mux_o_15_port, Z(14) => xor_mux_o_14_port, Z(13) => 
               xor_mux_o_13_port, Z(12) => xor_mux_o_12_port, Z(11) => 
               xor_mux_o_11_port, Z(10) => xor_mux_o_10_port, Z(9) => 
               xor_mux_o_9_port, Z(8) => xor_mux_o_8_port, Z(7) => 
               xor_mux_o_7_port, Z(6) => xor_mux_o_6_port, Z(5) => 
               xor_mux_o_5_port, Z(4) => xor_mux_o_4_port, Z(3) => 
               xor_mux_o_3_port, Z(2) => xor_mux_o_2_port, Z(1) => 
               xor_mux_o_1_port, Z(0) => xor_mux_o_0_port );
   B_8 : GTECH_BUF port map( A => N572, Z => N8);
   B_9 : GTECH_BUF port map( A => xor_sel, Z => N9);
   C1638_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 32 )
      port map(
         -- Connections to port 'DATA1'
         DATA(31) => temp_ram_31_port, DATA(30) => temp_ram_30_port, DATA(29) 
               => temp_ram_29_port, DATA(28) => temp_ram_28_port, DATA(27) => 
               temp_ram_27_port, DATA(26) => temp_ram_26_port, DATA(25) => 
               temp_ram_25_port, DATA(24) => temp_ram_24_port, DATA(23) => 
               temp_ram_23_port, DATA(22) => temp_ram_22_port, DATA(21) => 
               temp_ram_21_port, DATA(20) => temp_ram_20_port, DATA(19) => 
               temp_ram_19_port, DATA(18) => temp_ram_18_port, DATA(17) => 
               temp_ram_17_port, DATA(16) => temp_ram_16_port, DATA(15) => 
               temp_ram_15_port, DATA(14) => temp_ram_14_port, DATA(13) => 
               temp_ram_13_port, DATA(12) => temp_ram_12_port, DATA(11) => 
               temp_ram_11_port, DATA(10) => temp_ram_10_port, DATA(9) => 
               temp_ram_9_port, DATA(8) => temp_ram_8_port, DATA(7) => 
               temp_ram_7_port, DATA(6) => temp_ram_6_port, DATA(5) => 
               temp_ram_5_port, DATA(4) => temp_ram_4_port, DATA(3) => 
               temp_ram_3_port, DATA(2) => temp_ram_2_port, DATA(1) => 
               temp_ram_1_port, DATA(0) => temp_ram_0_port, 
         -- Connections to port 'DATA2'
         DATA(63) => temp_xor_out_31_port, DATA(62) => temp_xor_out_30_port, 
               DATA(61) => temp_xor_out_29_port, DATA(60) => 
               temp_xor_out_28_port, DATA(59) => temp_xor_out_27_port, DATA(58)
               => temp_xor_out_26_port, DATA(57) => temp_xor_out_25_port, 
               DATA(56) => temp_xor_out_24_port, DATA(55) => 
               temp_xor_out_23_port, DATA(54) => temp_xor_out_22_port, DATA(53)
               => temp_xor_out_21_port, DATA(52) => temp_xor_out_20_port, 
               DATA(51) => temp_xor_out_19_port, DATA(50) => 
               temp_xor_out_18_port, DATA(49) => temp_xor_out_17_port, DATA(48)
               => temp_xor_out_16_port, DATA(47) => temp_xor_out_15_port, 
               DATA(46) => temp_xor_out_14_port, DATA(45) => 
               temp_xor_out_13_port, DATA(44) => temp_xor_out_12_port, DATA(43)
               => temp_xor_out_11_port, DATA(42) => temp_xor_out_10_port, 
               DATA(41) => temp_xor_out_9_port, DATA(40) => temp_xor_out_8_port
               , DATA(39) => temp_xor_out_7_port, DATA(38) => 
               temp_xor_out_6_port, DATA(37) => temp_xor_out_5_port, DATA(36) 
               => temp_xor_out_4_port, DATA(35) => temp_xor_out_3_port, 
               DATA(34) => temp_xor_out_2_port, DATA(33) => temp_xor_out_1_port
               , DATA(32) => temp_xor_out_0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N10, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N11, 
         -- Connections to port 'Z'
         Z(31) => bdo_out_7_port, Z(30) => bdo_out_6_port, Z(29) => 
               bdo_out_5_port, Z(28) => bdo_out_4_port, Z(27) => bdo_out_3_port
               , Z(26) => bdo_out_2_port, Z(25) => bdo_out_1_port, Z(24) => 
               bdo_out_0_port, Z(23) => bdo_out_15_port, Z(22) => 
               bdo_out_14_port, Z(21) => bdo_out_13_port, Z(20) => 
               bdo_out_12_port, Z(19) => bdo_out_11_port, Z(18) => 
               bdo_out_10_port, Z(17) => bdo_out_9_port, Z(16) => 
               bdo_out_8_port, Z(15) => bdo_out_23_port, Z(14) => 
               bdo_out_22_port, Z(13) => bdo_out_21_port, Z(12) => 
               bdo_out_20_port, Z(11) => bdo_out_19_port, Z(10) => 
               bdo_out_18_port, Z(9) => bdo_out_17_port, Z(8) => 
               bdo_out_16_port, Z(7) => bdo_out_31_port, Z(6) => 
               bdo_out_30_port, Z(5) => bdo_out_29_port, Z(4) => 
               bdo_out_28_port, Z(3) => bdo_out_27_port, Z(2) => 
               bdo_out_26_port, Z(1) => bdo_out_25_port, Z(0) => 
               bdo_out_24_port );
   B_10 : GTECH_BUF port map( A => N571, Z => N10);
   B_11 : GTECH_BUF port map( A => extract_sel, Z => N11);
   C1639_cell : SELECT_OP
      generic map ( num_inputs => 4, input_width => 32 )
      port map(
         -- Connections to port 'DATA1'
         DATA(31) => plane_x_127_port, DATA(30) => plane_x_126_port, DATA(29) 
               => plane_x_125_port, DATA(28) => plane_x_124_port, DATA(27) => 
               plane_x_123_port, DATA(26) => plane_x_122_port, DATA(25) => 
               plane_x_121_port, DATA(24) => plane_x_120_port, DATA(23) => 
               plane_x_119_port, DATA(22) => plane_x_118_port, DATA(21) => 
               plane_x_117_port, DATA(20) => plane_x_116_port, DATA(19) => 
               plane_x_115_port, DATA(18) => plane_x_114_port, DATA(17) => 
               plane_x_113_port, DATA(16) => plane_x_112_port, DATA(15) => 
               plane_x_111_port, DATA(14) => plane_x_110_port, DATA(13) => 
               plane_x_109_port, DATA(12) => plane_x_108_port, DATA(11) => 
               plane_x_107_port, DATA(10) => plane_x_106_port, DATA(9) => 
               plane_x_105_port, DATA(8) => plane_x_104_port, DATA(7) => 
               plane_x_103_port, DATA(6) => plane_x_102_port, DATA(5) => 
               plane_x_101_port, DATA(4) => plane_x_100_port, DATA(3) => 
               plane_x_99_port, DATA(2) => plane_x_98_port, DATA(1) => 
               plane_x_97_port, DATA(0) => plane_x_96_port, 
         -- Connections to port 'DATA2'
         DATA(63) => plane_x_95_port, DATA(62) => plane_x_94_port, DATA(61) => 
               plane_x_93_port, DATA(60) => plane_x_92_port, DATA(59) => 
               plane_x_91_port, DATA(58) => plane_x_90_port, DATA(57) => 
               plane_x_89_port, DATA(56) => plane_x_88_port, DATA(55) => 
               plane_x_87_port, DATA(54) => plane_x_86_port, DATA(53) => 
               plane_x_85_port, DATA(52) => plane_x_84_port, DATA(51) => 
               plane_x_83_port, DATA(50) => plane_x_82_port, DATA(49) => 
               plane_x_81_port, DATA(48) => plane_x_80_port, DATA(47) => 
               plane_x_79_port, DATA(46) => plane_x_78_port, DATA(45) => 
               plane_x_77_port, DATA(44) => plane_x_76_port, DATA(43) => 
               plane_x_75_port, DATA(42) => plane_x_74_port, DATA(41) => 
               plane_x_73_port, DATA(40) => plane_x_72_port, DATA(39) => 
               plane_x_71_port, DATA(38) => plane_x_70_port, DATA(37) => 
               plane_x_69_port, DATA(36) => plane_x_68_port, DATA(35) => 
               plane_x_67_port, DATA(34) => plane_x_66_port, DATA(33) => 
               plane_x_65_port, DATA(32) => plane_x_64_port, 
         -- Connections to port 'DATA3'
         DATA(95) => plane_x_63_port, DATA(94) => plane_x_62_port, DATA(93) => 
               plane_x_61_port, DATA(92) => plane_x_60_port, DATA(91) => 
               plane_x_59_port, DATA(90) => plane_x_58_port, DATA(89) => 
               plane_x_57_port, DATA(88) => plane_x_56_port, DATA(87) => 
               plane_x_55_port, DATA(86) => plane_x_54_port, DATA(85) => 
               plane_x_53_port, DATA(84) => plane_x_52_port, DATA(83) => 
               plane_x_51_port, DATA(82) => plane_x_50_port, DATA(81) => 
               plane_x_49_port, DATA(80) => plane_x_48_port, DATA(79) => 
               plane_x_47_port, DATA(78) => plane_x_46_port, DATA(77) => 
               plane_x_45_port, DATA(76) => plane_x_44_port, DATA(75) => 
               plane_x_43_port, DATA(74) => plane_x_42_port, DATA(73) => 
               plane_x_41_port, DATA(72) => plane_x_40_port, DATA(71) => 
               plane_x_39_port, DATA(70) => plane_x_38_port, DATA(69) => 
               plane_x_37_port, DATA(68) => plane_x_36_port, DATA(67) => 
               plane_x_35_port, DATA(66) => plane_x_34_port, DATA(65) => 
               plane_x_33_port, DATA(64) => plane_x_32_port, 
         -- Connections to port 'DATA4'
         DATA(127) => plane_x_31_port, DATA(126) => plane_x_30_port, DATA(125) 
               => plane_x_29_port, DATA(124) => plane_x_28_port, DATA(123) => 
               plane_x_27_port, DATA(122) => plane_x_26_port, DATA(121) => 
               plane_x_25_port, DATA(120) => plane_x_24_port, DATA(119) => 
               plane_x_23_port, DATA(118) => plane_x_22_port, DATA(117) => 
               plane_x_21_port, DATA(116) => plane_x_20_port, DATA(115) => 
               plane_x_19_port, DATA(114) => plane_x_18_port, DATA(113) => 
               plane_x_17_port, DATA(112) => plane_x_16_port, DATA(111) => 
               plane_x_15_port, DATA(110) => plane_x_14_port, DATA(109) => 
               plane_x_13_port, DATA(108) => plane_x_12_port, DATA(107) => 
               plane_x_11_port, DATA(106) => plane_x_10_port, DATA(105) => 
               plane_x_9_port, DATA(104) => plane_x_8_port, DATA(103) => 
               plane_x_7_port, DATA(102) => plane_x_6_port, DATA(101) => 
               plane_x_5_port, DATA(100) => plane_x_4_port, DATA(99) => 
               plane_x_3_port, DATA(98) => plane_x_2_port, DATA(97) => 
               plane_x_1_port, DATA(96) => plane_x_0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N12, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N13, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N14, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N15, 
         -- Connections to port 'Z'
         Z(31) => temp_ram_31_port, Z(30) => temp_ram_30_port, Z(29) => 
               temp_ram_29_port, Z(28) => temp_ram_28_port, Z(27) => 
               temp_ram_27_port, Z(26) => temp_ram_26_port, Z(25) => 
               temp_ram_25_port, Z(24) => temp_ram_24_port, Z(23) => 
               temp_ram_23_port, Z(22) => temp_ram_22_port, Z(21) => 
               temp_ram_21_port, Z(20) => temp_ram_20_port, Z(19) => 
               temp_ram_19_port, Z(18) => temp_ram_18_port, Z(17) => 
               temp_ram_17_port, Z(16) => temp_ram_16_port, Z(15) => 
               temp_ram_15_port, Z(14) => temp_ram_14_port, Z(13) => 
               temp_ram_13_port, Z(12) => temp_ram_12_port, Z(11) => 
               temp_ram_11_port, Z(10) => temp_ram_10_port, Z(9) => 
               temp_ram_9_port, Z(8) => temp_ram_8_port, Z(7) => 
               temp_ram_7_port, Z(6) => temp_ram_6_port, Z(5) => 
               temp_ram_5_port, Z(4) => temp_ram_4_port, Z(3) => 
               temp_ram_3_port, Z(2) => temp_ram_2_port, Z(1) => 
               temp_ram_1_port, Z(0) => temp_ram_0_port );
   B_12 : GTECH_BUF port map( A => N172, Z => N12);
   B_13 : GTECH_BUF port map( A => N174, Z => N13);
   B_14 : GTECH_BUF port map( A => N176, Z => N14);
   B_15 : GTECH_BUF port map( A => N177, Z => N15);
   C1640_cell : SELECT_OP
      generic map ( num_inputs => 4, input_width => 24 )
      port map(
         -- Connections to port 'DATA1'
         DATA(23) => temp_ram_31_port, DATA(22) => temp_ram_30_port, DATA(21) 
               => temp_ram_29_port, DATA(20) => temp_ram_28_port, DATA(19) => 
               temp_ram_27_port, DATA(18) => temp_ram_26_port, DATA(17) => 
               temp_ram_25_port, DATA(16) => temp_ram_24_port, DATA(15) => 
               temp_ram_23_port, DATA(14) => temp_ram_22_port, DATA(13) => 
               temp_ram_21_port, DATA(12) => temp_ram_20_port, DATA(11) => 
               temp_ram_19_port, DATA(10) => temp_ram_18_port, DATA(9) => 
               temp_ram_17_port, DATA(8) => temp_ram_16_port, DATA(7) => 
               temp_ram_15_port, DATA(6) => temp_ram_14_port, DATA(5) => 
               temp_ram_13_port, DATA(4) => temp_ram_12_port, DATA(3) => 
               temp_ram_11_port, DATA(2) => temp_ram_10_port, DATA(1) => 
               temp_ram_9_port, DATA(0) => N178, 
         -- Connections to port 'DATA2'
         DATA(47) => temp_ram_31_port, DATA(46) => temp_ram_30_port, DATA(45) 
               => temp_ram_29_port, DATA(44) => temp_ram_28_port, DATA(43) => 
               temp_ram_27_port, DATA(42) => temp_ram_26_port, DATA(41) => 
               temp_ram_25_port, DATA(40) => temp_ram_24_port, DATA(39) => 
               temp_ram_23_port, DATA(38) => temp_ram_22_port, DATA(37) => 
               temp_ram_21_port, DATA(36) => temp_ram_20_port, DATA(35) => 
               temp_ram_19_port, DATA(34) => temp_ram_18_port, DATA(33) => 
               temp_ram_17_port, DATA(32) => N179, DATA(31) => bdi_key_23_port,
               DATA(30) => bdi_key_22_port, DATA(29) => bdi_key_21_port, 
               DATA(28) => bdi_key_20_port, DATA(27) => bdi_key_19_port, 
               DATA(26) => bdi_key_18_port, DATA(25) => bdi_key_17_port, 
               DATA(24) => bdi_key_16_port, 
         -- Connections to port 'DATA3'
         DATA(71) => temp_ram_31_port, DATA(70) => temp_ram_30_port, DATA(69) 
               => temp_ram_29_port, DATA(68) => temp_ram_28_port, DATA(67) => 
               temp_ram_27_port, DATA(66) => temp_ram_26_port, DATA(65) => 
               temp_ram_25_port, DATA(64) => N180, DATA(63) => bdi_key_15_port,
               DATA(62) => bdi_key_14_port, DATA(61) => bdi_key_13_port, 
               DATA(60) => bdi_key_12_port, DATA(59) => bdi_key_11_port, 
               DATA(58) => bdi_key_10_port, DATA(57) => bdi_key_9_port, 
               DATA(56) => bdi_key_8_port, DATA(55) => bdi_key_23_port, 
               DATA(54) => bdi_key_22_port, DATA(53) => bdi_key_21_port, 
               DATA(52) => bdi_key_20_port, DATA(51) => bdi_key_19_port, 
               DATA(50) => bdi_key_18_port, DATA(49) => bdi_key_17_port, 
               DATA(48) => bdi_key_16_port, 
         -- Connections to port 'DATA4'
         DATA(95) => bdi_key_7_port, DATA(94) => bdi_key_6_port, DATA(93) => 
               bdi_key_5_port, DATA(92) => bdi_key_4_port, DATA(91) => 
               bdi_key_3_port, DATA(90) => bdi_key_2_port, DATA(89) => 
               bdi_key_1_port, DATA(88) => bdi_key_0_port, DATA(87) => 
               bdi_key_15_port, DATA(86) => bdi_key_14_port, DATA(85) => 
               bdi_key_13_port, DATA(84) => bdi_key_12_port, DATA(83) => 
               bdi_key_11_port, DATA(82) => bdi_key_10_port, DATA(81) => 
               bdi_key_9_port, DATA(80) => bdi_key_8_port, DATA(79) => 
               bdi_key_23_port, DATA(78) => bdi_key_22_port, DATA(77) => 
               bdi_key_21_port, DATA(76) => bdi_key_20_port, DATA(75) => 
               bdi_key_19_port, DATA(74) => bdi_key_18_port, DATA(73) => 
               bdi_key_17_port, DATA(72) => bdi_key_16_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N4, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N5, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N6, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N7, 
         -- Connections to port 'Z'
         Z(23) => decrypt_mux_31_port, Z(22) => decrypt_mux_30_port, Z(21) => 
               decrypt_mux_29_port, Z(20) => decrypt_mux_28_port, Z(19) => 
               decrypt_mux_27_port, Z(18) => decrypt_mux_26_port, Z(17) => 
               decrypt_mux_25_port, Z(16) => decrypt_mux_24_port, Z(15) => 
               decrypt_mux_23_port, Z(14) => decrypt_mux_22_port, Z(13) => 
               decrypt_mux_21_port, Z(12) => decrypt_mux_20_port, Z(11) => 
               decrypt_mux_19_port, Z(10) => decrypt_mux_18_port, Z(9) => 
               decrypt_mux_17_port, Z(8) => decrypt_mux_16_port, Z(7) => 
               decrypt_mux_15_port, Z(6) => decrypt_mux_14_port, Z(5) => 
               decrypt_mux_13_port, Z(4) => decrypt_mux_12_port, Z(3) => 
               decrypt_mux_11_port, Z(2) => decrypt_mux_10_port, Z(1) => 
               decrypt_mux_9_port, Z(0) => decrypt_mux_8_port );
   C1641_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 32 )
      port map(
         -- Connections to port 'DATA1'
         DATA(31) => temp_xor_out_31_port, DATA(30) => temp_xor_out_30_port, 
               DATA(29) => temp_xor_out_29_port, DATA(28) => 
               temp_xor_out_28_port, DATA(27) => temp_xor_out_27_port, DATA(26)
               => temp_xor_out_26_port, DATA(25) => temp_xor_out_25_port, 
               DATA(24) => temp_xor_out_24_port, DATA(23) => 
               temp_xor_out_23_port, DATA(22) => temp_xor_out_22_port, DATA(21)
               => temp_xor_out_21_port, DATA(20) => temp_xor_out_20_port, 
               DATA(19) => temp_xor_out_19_port, DATA(18) => 
               temp_xor_out_18_port, DATA(17) => temp_xor_out_17_port, DATA(16)
               => temp_xor_out_16_port, DATA(15) => temp_xor_out_15_port, 
               DATA(14) => temp_xor_out_14_port, DATA(13) => 
               temp_xor_out_13_port, DATA(12) => temp_xor_out_12_port, DATA(11)
               => temp_xor_out_11_port, DATA(10) => temp_xor_out_10_port, 
               DATA(9) => temp_xor_out_9_port, DATA(8) => temp_xor_out_8_port, 
               DATA(7) => temp_xor_out_7_port, DATA(6) => temp_xor_out_6_port, 
               DATA(5) => temp_xor_out_5_port, DATA(4) => temp_xor_out_4_port, 
               DATA(3) => temp_xor_out_3_port, DATA(2) => temp_xor_out_2_port, 
               DATA(1) => temp_xor_out_1_port, DATA(0) => temp_xor_out_0_port, 
         -- Connections to port 'DATA2'
         DATA(63) => decrypt_mux_31_port, DATA(62) => decrypt_mux_30_port, 
               DATA(61) => decrypt_mux_29_port, DATA(60) => decrypt_mux_28_port
               , DATA(59) => decrypt_mux_27_port, DATA(58) => 
               decrypt_mux_26_port, DATA(57) => decrypt_mux_25_port, DATA(56) 
               => decrypt_mux_24_port, DATA(55) => decrypt_mux_23_port, 
               DATA(54) => decrypt_mux_22_port, DATA(53) => decrypt_mux_21_port
               , DATA(52) => decrypt_mux_20_port, DATA(51) => 
               decrypt_mux_19_port, DATA(50) => decrypt_mux_18_port, DATA(49) 
               => decrypt_mux_17_port, DATA(48) => decrypt_mux_16_port, 
               DATA(47) => decrypt_mux_15_port, DATA(46) => decrypt_mux_14_port
               , DATA(45) => decrypt_mux_13_port, DATA(44) => 
               decrypt_mux_12_port, DATA(43) => decrypt_mux_11_port, DATA(42) 
               => decrypt_mux_10_port, DATA(41) => decrypt_mux_9_port, DATA(40)
               => decrypt_mux_8_port, DATA(39) => bdi_key_31_port, DATA(38) => 
               bdi_key_30_port, DATA(37) => bdi_key_29_port, DATA(36) => 
               bdi_key_28_port, DATA(35) => bdi_key_27_port, DATA(34) => 
               bdi_key_26_port, DATA(33) => bdi_key_25_port, DATA(32) => 
               bdi_key_24_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N16, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N17, 
         -- Connections to port 'Z'
         Z(31) => temp_cyc_state_31_port, Z(30) => temp_cyc_state_30_port, 
               Z(29) => temp_cyc_state_29_port, Z(28) => temp_cyc_state_28_port
               , Z(27) => temp_cyc_state_27_port, Z(26) => 
               temp_cyc_state_26_port, Z(25) => temp_cyc_state_25_port, Z(24) 
               => temp_cyc_state_24_port, Z(23) => temp_cyc_state_23_port, 
               Z(22) => temp_cyc_state_22_port, Z(21) => temp_cyc_state_21_port
               , Z(20) => temp_cyc_state_20_port, Z(19) => 
               temp_cyc_state_19_port, Z(18) => temp_cyc_state_18_port, Z(17) 
               => temp_cyc_state_17_port, Z(16) => temp_cyc_state_16_port, 
               Z(15) => temp_cyc_state_15_port, Z(14) => temp_cyc_state_14_port
               , Z(13) => temp_cyc_state_13_port, Z(12) => 
               temp_cyc_state_12_port, Z(11) => temp_cyc_state_11_port, Z(10) 
               => temp_cyc_state_10_port, Z(9) => temp_cyc_state_9_port, Z(8) 
               => temp_cyc_state_8_port, Z(7) => temp_cyc_state_7_port, Z(6) =>
               temp_cyc_state_6_port, Z(5) => temp_cyc_state_5_port, Z(4) => 
               temp_cyc_state_4_port, Z(3) => temp_cyc_state_3_port, Z(2) => 
               temp_cyc_state_2_port, Z(1) => temp_cyc_state_1_port, Z(0) => 
               temp_cyc_state_0_port );
   B_16 : GTECH_BUF port map( A => N573, Z => N16);
   B_17 : GTECH_BUF port map( A => cyc_state_update_sel, Z => N17);
   C1642_cell : SELECT_OP
      generic map ( num_inputs => 4, input_width => 128 )
      port map(
         -- Connections to port 'DATA1'
         DATA(127) => temp_cyc_state_31_port, DATA(126) => 
               temp_cyc_state_30_port, DATA(125) => temp_cyc_state_29_port, 
               DATA(124) => temp_cyc_state_28_port, DATA(123) => 
               temp_cyc_state_27_port, DATA(122) => temp_cyc_state_26_port, 
               DATA(121) => temp_cyc_state_25_port, DATA(120) => 
               temp_cyc_state_24_port, DATA(119) => temp_cyc_state_23_port, 
               DATA(118) => temp_cyc_state_22_port, DATA(117) => 
               temp_cyc_state_21_port, DATA(116) => temp_cyc_state_20_port, 
               DATA(115) => temp_cyc_state_19_port, DATA(114) => 
               temp_cyc_state_18_port, DATA(113) => temp_cyc_state_17_port, 
               DATA(112) => temp_cyc_state_16_port, DATA(111) => 
               temp_cyc_state_15_port, DATA(110) => temp_cyc_state_14_port, 
               DATA(109) => temp_cyc_state_13_port, DATA(108) => 
               temp_cyc_state_12_port, DATA(107) => temp_cyc_state_11_port, 
               DATA(106) => temp_cyc_state_10_port, DATA(105) => 
               temp_cyc_state_9_port, DATA(104) => temp_cyc_state_8_port, 
               DATA(103) => temp_cyc_state_7_port, DATA(102) => 
               temp_cyc_state_6_port, DATA(101) => temp_cyc_state_5_port, 
               DATA(100) => temp_cyc_state_4_port, DATA(99) => 
               temp_cyc_state_3_port, DATA(98) => temp_cyc_state_2_port, 
               DATA(97) => temp_cyc_state_1_port, DATA(96) => 
               temp_cyc_state_0_port, DATA(95) => plane_x_95_port, DATA(94) => 
               plane_x_94_port, DATA(93) => plane_x_93_port, DATA(92) => 
               plane_x_92_port, DATA(91) => plane_x_91_port, DATA(90) => 
               plane_x_90_port, DATA(89) => plane_x_89_port, DATA(88) => 
               plane_x_88_port, DATA(87) => plane_x_87_port, DATA(86) => 
               plane_x_86_port, DATA(85) => plane_x_85_port, DATA(84) => 
               plane_x_84_port, DATA(83) => plane_x_83_port, DATA(82) => 
               plane_x_82_port, DATA(81) => plane_x_81_port, DATA(80) => 
               plane_x_80_port, DATA(79) => plane_x_79_port, DATA(78) => 
               plane_x_78_port, DATA(77) => plane_x_77_port, DATA(76) => 
               plane_x_76_port, DATA(75) => plane_x_75_port, DATA(74) => 
               plane_x_74_port, DATA(73) => plane_x_73_port, DATA(72) => 
               plane_x_72_port, DATA(71) => plane_x_71_port, DATA(70) => 
               plane_x_70_port, DATA(69) => plane_x_69_port, DATA(68) => 
               plane_x_68_port, DATA(67) => plane_x_67_port, DATA(66) => 
               plane_x_66_port, DATA(65) => plane_x_65_port, DATA(64) => 
               plane_x_64_port, DATA(63) => plane_x_63_port, DATA(62) => 
               plane_x_62_port, DATA(61) => plane_x_61_port, DATA(60) => 
               plane_x_60_port, DATA(59) => plane_x_59_port, DATA(58) => 
               plane_x_58_port, DATA(57) => plane_x_57_port, DATA(56) => 
               plane_x_56_port, DATA(55) => plane_x_55_port, DATA(54) => 
               plane_x_54_port, DATA(53) => plane_x_53_port, DATA(52) => 
               plane_x_52_port, DATA(51) => plane_x_51_port, DATA(50) => 
               plane_x_50_port, DATA(49) => plane_x_49_port, DATA(48) => 
               plane_x_48_port, DATA(47) => plane_x_47_port, DATA(46) => 
               plane_x_46_port, DATA(45) => plane_x_45_port, DATA(44) => 
               plane_x_44_port, DATA(43) => plane_x_43_port, DATA(42) => 
               plane_x_42_port, DATA(41) => plane_x_41_port, DATA(40) => 
               plane_x_40_port, DATA(39) => plane_x_39_port, DATA(38) => 
               plane_x_38_port, DATA(37) => plane_x_37_port, DATA(36) => 
               plane_x_36_port, DATA(35) => plane_x_35_port, DATA(34) => 
               plane_x_34_port, DATA(33) => plane_x_33_port, DATA(32) => 
               plane_x_32_port, DATA(31) => plane_x_31_port, DATA(30) => 
               plane_x_30_port, DATA(29) => plane_x_29_port, DATA(28) => 
               plane_x_28_port, DATA(27) => plane_x_27_port, DATA(26) => 
               plane_x_26_port, DATA(25) => plane_x_25_port, DATA(24) => 
               plane_x_24_port, DATA(23) => plane_x_23_port, DATA(22) => 
               plane_x_22_port, DATA(21) => plane_x_21_port, DATA(20) => 
               plane_x_20_port, DATA(19) => plane_x_19_port, DATA(18) => 
               plane_x_18_port, DATA(17) => plane_x_17_port, DATA(16) => 
               plane_x_16_port, DATA(15) => plane_x_15_port, DATA(14) => 
               plane_x_14_port, DATA(13) => plane_x_13_port, DATA(12) => 
               plane_x_12_port, DATA(11) => plane_x_11_port, DATA(10) => 
               plane_x_10_port, DATA(9) => plane_x_9_port, DATA(8) => 
               plane_x_8_port, DATA(7) => plane_x_7_port, DATA(6) => 
               plane_x_6_port, DATA(5) => plane_x_5_port, DATA(4) => 
               plane_x_4_port, DATA(3) => plane_x_3_port, DATA(2) => 
               plane_x_2_port, DATA(1) => plane_x_1_port, DATA(0) => 
               plane_x_0_port, 
         -- Connections to port 'DATA2'
         DATA(255) => plane_x_127_port, DATA(254) => plane_x_126_port, 
               DATA(253) => plane_x_125_port, DATA(252) => plane_x_124_port, 
               DATA(251) => plane_x_123_port, DATA(250) => plane_x_122_port, 
               DATA(249) => plane_x_121_port, DATA(248) => plane_x_120_port, 
               DATA(247) => plane_x_119_port, DATA(246) => plane_x_118_port, 
               DATA(245) => plane_x_117_port, DATA(244) => plane_x_116_port, 
               DATA(243) => plane_x_115_port, DATA(242) => plane_x_114_port, 
               DATA(241) => plane_x_113_port, DATA(240) => plane_x_112_port, 
               DATA(239) => plane_x_111_port, DATA(238) => plane_x_110_port, 
               DATA(237) => plane_x_109_port, DATA(236) => plane_x_108_port, 
               DATA(235) => plane_x_107_port, DATA(234) => plane_x_106_port, 
               DATA(233) => plane_x_105_port, DATA(232) => plane_x_104_port, 
               DATA(231) => plane_x_103_port, DATA(230) => plane_x_102_port, 
               DATA(229) => plane_x_101_port, DATA(228) => plane_x_100_port, 
               DATA(227) => plane_x_99_port, DATA(226) => plane_x_98_port, 
               DATA(225) => plane_x_97_port, DATA(224) => plane_x_96_port, 
               DATA(223) => temp_cyc_state_31_port, DATA(222) => 
               temp_cyc_state_30_port, DATA(221) => temp_cyc_state_29_port, 
               DATA(220) => temp_cyc_state_28_port, DATA(219) => 
               temp_cyc_state_27_port, DATA(218) => temp_cyc_state_26_port, 
               DATA(217) => temp_cyc_state_25_port, DATA(216) => 
               temp_cyc_state_24_port, DATA(215) => temp_cyc_state_23_port, 
               DATA(214) => temp_cyc_state_22_port, DATA(213) => 
               temp_cyc_state_21_port, DATA(212) => temp_cyc_state_20_port, 
               DATA(211) => temp_cyc_state_19_port, DATA(210) => 
               temp_cyc_state_18_port, DATA(209) => temp_cyc_state_17_port, 
               DATA(208) => temp_cyc_state_16_port, DATA(207) => 
               temp_cyc_state_15_port, DATA(206) => temp_cyc_state_14_port, 
               DATA(205) => temp_cyc_state_13_port, DATA(204) => 
               temp_cyc_state_12_port, DATA(203) => temp_cyc_state_11_port, 
               DATA(202) => temp_cyc_state_10_port, DATA(201) => 
               temp_cyc_state_9_port, DATA(200) => temp_cyc_state_8_port, 
               DATA(199) => temp_cyc_state_7_port, DATA(198) => 
               temp_cyc_state_6_port, DATA(197) => temp_cyc_state_5_port, 
               DATA(196) => temp_cyc_state_4_port, DATA(195) => 
               temp_cyc_state_3_port, DATA(194) => temp_cyc_state_2_port, 
               DATA(193) => temp_cyc_state_1_port, DATA(192) => 
               temp_cyc_state_0_port, DATA(191) => plane_x_63_port, DATA(190) 
               => plane_x_62_port, DATA(189) => plane_x_61_port, DATA(188) => 
               plane_x_60_port, DATA(187) => plane_x_59_port, DATA(186) => 
               plane_x_58_port, DATA(185) => plane_x_57_port, DATA(184) => 
               plane_x_56_port, DATA(183) => plane_x_55_port, DATA(182) => 
               plane_x_54_port, DATA(181) => plane_x_53_port, DATA(180) => 
               plane_x_52_port, DATA(179) => plane_x_51_port, DATA(178) => 
               plane_x_50_port, DATA(177) => plane_x_49_port, DATA(176) => 
               plane_x_48_port, DATA(175) => plane_x_47_port, DATA(174) => 
               plane_x_46_port, DATA(173) => plane_x_45_port, DATA(172) => 
               plane_x_44_port, DATA(171) => plane_x_43_port, DATA(170) => 
               plane_x_42_port, DATA(169) => plane_x_41_port, DATA(168) => 
               plane_x_40_port, DATA(167) => plane_x_39_port, DATA(166) => 
               plane_x_38_port, DATA(165) => plane_x_37_port, DATA(164) => 
               plane_x_36_port, DATA(163) => plane_x_35_port, DATA(162) => 
               plane_x_34_port, DATA(161) => plane_x_33_port, DATA(160) => 
               plane_x_32_port, DATA(159) => plane_x_31_port, DATA(158) => 
               plane_x_30_port, DATA(157) => plane_x_29_port, DATA(156) => 
               plane_x_28_port, DATA(155) => plane_x_27_port, DATA(154) => 
               plane_x_26_port, DATA(153) => plane_x_25_port, DATA(152) => 
               plane_x_24_port, DATA(151) => plane_x_23_port, DATA(150) => 
               plane_x_22_port, DATA(149) => plane_x_21_port, DATA(148) => 
               plane_x_20_port, DATA(147) => plane_x_19_port, DATA(146) => 
               plane_x_18_port, DATA(145) => plane_x_17_port, DATA(144) => 
               plane_x_16_port, DATA(143) => plane_x_15_port, DATA(142) => 
               plane_x_14_port, DATA(141) => plane_x_13_port, DATA(140) => 
               plane_x_12_port, DATA(139) => plane_x_11_port, DATA(138) => 
               plane_x_10_port, DATA(137) => plane_x_9_port, DATA(136) => 
               plane_x_8_port, DATA(135) => plane_x_7_port, DATA(134) => 
               plane_x_6_port, DATA(133) => plane_x_5_port, DATA(132) => 
               plane_x_4_port, DATA(131) => plane_x_3_port, DATA(130) => 
               plane_x_2_port, DATA(129) => plane_x_1_port, DATA(128) => 
               plane_x_0_port, 
         -- Connections to port 'DATA3'
         DATA(383) => plane_x_127_port, DATA(382) => plane_x_126_port, 
               DATA(381) => plane_x_125_port, DATA(380) => plane_x_124_port, 
               DATA(379) => plane_x_123_port, DATA(378) => plane_x_122_port, 
               DATA(377) => plane_x_121_port, DATA(376) => plane_x_120_port, 
               DATA(375) => plane_x_119_port, DATA(374) => plane_x_118_port, 
               DATA(373) => plane_x_117_port, DATA(372) => plane_x_116_port, 
               DATA(371) => plane_x_115_port, DATA(370) => plane_x_114_port, 
               DATA(369) => plane_x_113_port, DATA(368) => plane_x_112_port, 
               DATA(367) => plane_x_111_port, DATA(366) => plane_x_110_port, 
               DATA(365) => plane_x_109_port, DATA(364) => plane_x_108_port, 
               DATA(363) => plane_x_107_port, DATA(362) => plane_x_106_port, 
               DATA(361) => plane_x_105_port, DATA(360) => plane_x_104_port, 
               DATA(359) => plane_x_103_port, DATA(358) => plane_x_102_port, 
               DATA(357) => plane_x_101_port, DATA(356) => plane_x_100_port, 
               DATA(355) => plane_x_99_port, DATA(354) => plane_x_98_port, 
               DATA(353) => plane_x_97_port, DATA(352) => plane_x_96_port, 
               DATA(351) => plane_x_95_port, DATA(350) => plane_x_94_port, 
               DATA(349) => plane_x_93_port, DATA(348) => plane_x_92_port, 
               DATA(347) => plane_x_91_port, DATA(346) => plane_x_90_port, 
               DATA(345) => plane_x_89_port, DATA(344) => plane_x_88_port, 
               DATA(343) => plane_x_87_port, DATA(342) => plane_x_86_port, 
               DATA(341) => plane_x_85_port, DATA(340) => plane_x_84_port, 
               DATA(339) => plane_x_83_port, DATA(338) => plane_x_82_port, 
               DATA(337) => plane_x_81_port, DATA(336) => plane_x_80_port, 
               DATA(335) => plane_x_79_port, DATA(334) => plane_x_78_port, 
               DATA(333) => plane_x_77_port, DATA(332) => plane_x_76_port, 
               DATA(331) => plane_x_75_port, DATA(330) => plane_x_74_port, 
               DATA(329) => plane_x_73_port, DATA(328) => plane_x_72_port, 
               DATA(327) => plane_x_71_port, DATA(326) => plane_x_70_port, 
               DATA(325) => plane_x_69_port, DATA(324) => plane_x_68_port, 
               DATA(323) => plane_x_67_port, DATA(322) => plane_x_66_port, 
               DATA(321) => plane_x_65_port, DATA(320) => plane_x_64_port, 
               DATA(319) => temp_cyc_state_31_port, DATA(318) => 
               temp_cyc_state_30_port, DATA(317) => temp_cyc_state_29_port, 
               DATA(316) => temp_cyc_state_28_port, DATA(315) => 
               temp_cyc_state_27_port, DATA(314) => temp_cyc_state_26_port, 
               DATA(313) => temp_cyc_state_25_port, DATA(312) => 
               temp_cyc_state_24_port, DATA(311) => temp_cyc_state_23_port, 
               DATA(310) => temp_cyc_state_22_port, DATA(309) => 
               temp_cyc_state_21_port, DATA(308) => temp_cyc_state_20_port, 
               DATA(307) => temp_cyc_state_19_port, DATA(306) => 
               temp_cyc_state_18_port, DATA(305) => temp_cyc_state_17_port, 
               DATA(304) => temp_cyc_state_16_port, DATA(303) => 
               temp_cyc_state_15_port, DATA(302) => temp_cyc_state_14_port, 
               DATA(301) => temp_cyc_state_13_port, DATA(300) => 
               temp_cyc_state_12_port, DATA(299) => temp_cyc_state_11_port, 
               DATA(298) => temp_cyc_state_10_port, DATA(297) => 
               temp_cyc_state_9_port, DATA(296) => temp_cyc_state_8_port, 
               DATA(295) => temp_cyc_state_7_port, DATA(294) => 
               temp_cyc_state_6_port, DATA(293) => temp_cyc_state_5_port, 
               DATA(292) => temp_cyc_state_4_port, DATA(291) => 
               temp_cyc_state_3_port, DATA(290) => temp_cyc_state_2_port, 
               DATA(289) => temp_cyc_state_1_port, DATA(288) => 
               temp_cyc_state_0_port, DATA(287) => plane_x_31_port, DATA(286) 
               => plane_x_30_port, DATA(285) => plane_x_29_port, DATA(284) => 
               plane_x_28_port, DATA(283) => plane_x_27_port, DATA(282) => 
               plane_x_26_port, DATA(281) => plane_x_25_port, DATA(280) => 
               plane_x_24_port, DATA(279) => plane_x_23_port, DATA(278) => 
               plane_x_22_port, DATA(277) => plane_x_21_port, DATA(276) => 
               plane_x_20_port, DATA(275) => plane_x_19_port, DATA(274) => 
               plane_x_18_port, DATA(273) => plane_x_17_port, DATA(272) => 
               plane_x_16_port, DATA(271) => plane_x_15_port, DATA(270) => 
               plane_x_14_port, DATA(269) => plane_x_13_port, DATA(268) => 
               plane_x_12_port, DATA(267) => plane_x_11_port, DATA(266) => 
               plane_x_10_port, DATA(265) => plane_x_9_port, DATA(264) => 
               plane_x_8_port, DATA(263) => plane_x_7_port, DATA(262) => 
               plane_x_6_port, DATA(261) => plane_x_5_port, DATA(260) => 
               plane_x_4_port, DATA(259) => plane_x_3_port, DATA(258) => 
               plane_x_2_port, DATA(257) => plane_x_1_port, DATA(256) => 
               plane_x_0_port, 
         -- Connections to port 'DATA4'
         DATA(511) => plane_x_127_port, DATA(510) => plane_x_126_port, 
               DATA(509) => plane_x_125_port, DATA(508) => plane_x_124_port, 
               DATA(507) => plane_x_123_port, DATA(506) => plane_x_122_port, 
               DATA(505) => plane_x_121_port, DATA(504) => plane_x_120_port, 
               DATA(503) => plane_x_119_port, DATA(502) => plane_x_118_port, 
               DATA(501) => plane_x_117_port, DATA(500) => plane_x_116_port, 
               DATA(499) => plane_x_115_port, DATA(498) => plane_x_114_port, 
               DATA(497) => plane_x_113_port, DATA(496) => plane_x_112_port, 
               DATA(495) => plane_x_111_port, DATA(494) => plane_x_110_port, 
               DATA(493) => plane_x_109_port, DATA(492) => plane_x_108_port, 
               DATA(491) => plane_x_107_port, DATA(490) => plane_x_106_port, 
               DATA(489) => plane_x_105_port, DATA(488) => plane_x_104_port, 
               DATA(487) => plane_x_103_port, DATA(486) => plane_x_102_port, 
               DATA(485) => plane_x_101_port, DATA(484) => plane_x_100_port, 
               DATA(483) => plane_x_99_port, DATA(482) => plane_x_98_port, 
               DATA(481) => plane_x_97_port, DATA(480) => plane_x_96_port, 
               DATA(479) => plane_x_95_port, DATA(478) => plane_x_94_port, 
               DATA(477) => plane_x_93_port, DATA(476) => plane_x_92_port, 
               DATA(475) => plane_x_91_port, DATA(474) => plane_x_90_port, 
               DATA(473) => plane_x_89_port, DATA(472) => plane_x_88_port, 
               DATA(471) => plane_x_87_port, DATA(470) => plane_x_86_port, 
               DATA(469) => plane_x_85_port, DATA(468) => plane_x_84_port, 
               DATA(467) => plane_x_83_port, DATA(466) => plane_x_82_port, 
               DATA(465) => plane_x_81_port, DATA(464) => plane_x_80_port, 
               DATA(463) => plane_x_79_port, DATA(462) => plane_x_78_port, 
               DATA(461) => plane_x_77_port, DATA(460) => plane_x_76_port, 
               DATA(459) => plane_x_75_port, DATA(458) => plane_x_74_port, 
               DATA(457) => plane_x_73_port, DATA(456) => plane_x_72_port, 
               DATA(455) => plane_x_71_port, DATA(454) => plane_x_70_port, 
               DATA(453) => plane_x_69_port, DATA(452) => plane_x_68_port, 
               DATA(451) => plane_x_67_port, DATA(450) => plane_x_66_port, 
               DATA(449) => plane_x_65_port, DATA(448) => plane_x_64_port, 
               DATA(447) => plane_x_63_port, DATA(446) => plane_x_62_port, 
               DATA(445) => plane_x_61_port, DATA(444) => plane_x_60_port, 
               DATA(443) => plane_x_59_port, DATA(442) => plane_x_58_port, 
               DATA(441) => plane_x_57_port, DATA(440) => plane_x_56_port, 
               DATA(439) => plane_x_55_port, DATA(438) => plane_x_54_port, 
               DATA(437) => plane_x_53_port, DATA(436) => plane_x_52_port, 
               DATA(435) => plane_x_51_port, DATA(434) => plane_x_50_port, 
               DATA(433) => plane_x_49_port, DATA(432) => plane_x_48_port, 
               DATA(431) => plane_x_47_port, DATA(430) => plane_x_46_port, 
               DATA(429) => plane_x_45_port, DATA(428) => plane_x_44_port, 
               DATA(427) => plane_x_43_port, DATA(426) => plane_x_42_port, 
               DATA(425) => plane_x_41_port, DATA(424) => plane_x_40_port, 
               DATA(423) => plane_x_39_port, DATA(422) => plane_x_38_port, 
               DATA(421) => plane_x_37_port, DATA(420) => plane_x_36_port, 
               DATA(419) => plane_x_35_port, DATA(418) => plane_x_34_port, 
               DATA(417) => plane_x_33_port, DATA(416) => plane_x_32_port, 
               DATA(415) => temp_cyc_state_31_port, DATA(414) => 
               temp_cyc_state_30_port, DATA(413) => temp_cyc_state_29_port, 
               DATA(412) => temp_cyc_state_28_port, DATA(411) => 
               temp_cyc_state_27_port, DATA(410) => temp_cyc_state_26_port, 
               DATA(409) => temp_cyc_state_25_port, DATA(408) => 
               temp_cyc_state_24_port, DATA(407) => temp_cyc_state_23_port, 
               DATA(406) => temp_cyc_state_22_port, DATA(405) => 
               temp_cyc_state_21_port, DATA(404) => temp_cyc_state_20_port, 
               DATA(403) => temp_cyc_state_19_port, DATA(402) => 
               temp_cyc_state_18_port, DATA(401) => temp_cyc_state_17_port, 
               DATA(400) => temp_cyc_state_16_port, DATA(399) => 
               temp_cyc_state_15_port, DATA(398) => temp_cyc_state_14_port, 
               DATA(397) => temp_cyc_state_13_port, DATA(396) => 
               temp_cyc_state_12_port, DATA(395) => temp_cyc_state_11_port, 
               DATA(394) => temp_cyc_state_10_port, DATA(393) => 
               temp_cyc_state_9_port, DATA(392) => temp_cyc_state_8_port, 
               DATA(391) => temp_cyc_state_7_port, DATA(390) => 
               temp_cyc_state_6_port, DATA(389) => temp_cyc_state_5_port, 
               DATA(388) => temp_cyc_state_4_port, DATA(387) => 
               temp_cyc_state_3_port, DATA(386) => temp_cyc_state_2_port, 
               DATA(385) => temp_cyc_state_1_port, DATA(384) => 
               temp_cyc_state_0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N12, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N13, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N14, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N15, 
         -- Connections to port 'Z'
         Z(127) => cyc_state_update_127_port, Z(126) => 
               cyc_state_update_126_port, Z(125) => cyc_state_update_125_port, 
               Z(124) => cyc_state_update_124_port, Z(123) => 
               cyc_state_update_123_port, Z(122) => cyc_state_update_122_port, 
               Z(121) => cyc_state_update_121_port, Z(120) => 
               cyc_state_update_120_port, Z(119) => cyc_state_update_119_port, 
               Z(118) => cyc_state_update_118_port, Z(117) => 
               cyc_state_update_117_port, Z(116) => cyc_state_update_116_port, 
               Z(115) => cyc_state_update_115_port, Z(114) => 
               cyc_state_update_114_port, Z(113) => cyc_state_update_113_port, 
               Z(112) => cyc_state_update_112_port, Z(111) => 
               cyc_state_update_111_port, Z(110) => cyc_state_update_110_port, 
               Z(109) => cyc_state_update_109_port, Z(108) => 
               cyc_state_update_108_port, Z(107) => cyc_state_update_107_port, 
               Z(106) => cyc_state_update_106_port, Z(105) => 
               cyc_state_update_105_port, Z(104) => cyc_state_update_104_port, 
               Z(103) => cyc_state_update_103_port, Z(102) => 
               cyc_state_update_102_port, Z(101) => cyc_state_update_101_port, 
               Z(100) => cyc_state_update_100_port, Z(99) => 
               cyc_state_update_99_port, Z(98) => cyc_state_update_98_port, 
               Z(97) => cyc_state_update_97_port, Z(96) => 
               cyc_state_update_96_port, Z(95) => cyc_state_update_95_port, 
               Z(94) => cyc_state_update_94_port, Z(93) => 
               cyc_state_update_93_port, Z(92) => cyc_state_update_92_port, 
               Z(91) => cyc_state_update_91_port, Z(90) => 
               cyc_state_update_90_port, Z(89) => cyc_state_update_89_port, 
               Z(88) => cyc_state_update_88_port, Z(87) => 
               cyc_state_update_87_port, Z(86) => cyc_state_update_86_port, 
               Z(85) => cyc_state_update_85_port, Z(84) => 
               cyc_state_update_84_port, Z(83) => cyc_state_update_83_port, 
               Z(82) => cyc_state_update_82_port, Z(81) => 
               cyc_state_update_81_port, Z(80) => cyc_state_update_80_port, 
               Z(79) => cyc_state_update_79_port, Z(78) => 
               cyc_state_update_78_port, Z(77) => cyc_state_update_77_port, 
               Z(76) => cyc_state_update_76_port, Z(75) => 
               cyc_state_update_75_port, Z(74) => cyc_state_update_74_port, 
               Z(73) => cyc_state_update_73_port, Z(72) => 
               cyc_state_update_72_port, Z(71) => cyc_state_update_71_port, 
               Z(70) => cyc_state_update_70_port, Z(69) => 
               cyc_state_update_69_port, Z(68) => cyc_state_update_68_port, 
               Z(67) => cyc_state_update_67_port, Z(66) => 
               cyc_state_update_66_port, Z(65) => cyc_state_update_65_port, 
               Z(64) => cyc_state_update_64_port, Z(63) => 
               cyc_state_update_63_port, Z(62) => cyc_state_update_62_port, 
               Z(61) => cyc_state_update_61_port, Z(60) => 
               cyc_state_update_60_port, Z(59) => cyc_state_update_59_port, 
               Z(58) => cyc_state_update_58_port, Z(57) => 
               cyc_state_update_57_port, Z(56) => cyc_state_update_56_port, 
               Z(55) => cyc_state_update_55_port, Z(54) => 
               cyc_state_update_54_port, Z(53) => cyc_state_update_53_port, 
               Z(52) => cyc_state_update_52_port, Z(51) => 
               cyc_state_update_51_port, Z(50) => cyc_state_update_50_port, 
               Z(49) => cyc_state_update_49_port, Z(48) => 
               cyc_state_update_48_port, Z(47) => cyc_state_update_47_port, 
               Z(46) => cyc_state_update_46_port, Z(45) => 
               cyc_state_update_45_port, Z(44) => cyc_state_update_44_port, 
               Z(43) => cyc_state_update_43_port, Z(42) => 
               cyc_state_update_42_port, Z(41) => cyc_state_update_41_port, 
               Z(40) => cyc_state_update_40_port, Z(39) => 
               cyc_state_update_39_port, Z(38) => cyc_state_update_38_port, 
               Z(37) => cyc_state_update_37_port, Z(36) => 
               cyc_state_update_36_port, Z(35) => cyc_state_update_35_port, 
               Z(34) => cyc_state_update_34_port, Z(33) => 
               cyc_state_update_33_port, Z(32) => cyc_state_update_32_port, 
               Z(31) => cyc_state_update_31_port, Z(30) => 
               cyc_state_update_30_port, Z(29) => cyc_state_update_29_port, 
               Z(28) => cyc_state_update_28_port, Z(27) => 
               cyc_state_update_27_port, Z(26) => cyc_state_update_26_port, 
               Z(25) => cyc_state_update_25_port, Z(24) => 
               cyc_state_update_24_port, Z(23) => cyc_state_update_23_port, 
               Z(22) => cyc_state_update_22_port, Z(21) => 
               cyc_state_update_21_port, Z(20) => cyc_state_update_20_port, 
               Z(19) => cyc_state_update_19_port, Z(18) => 
               cyc_state_update_18_port, Z(17) => cyc_state_update_17_port, 
               Z(16) => cyc_state_update_16_port, Z(15) => 
               cyc_state_update_15_port, Z(14) => cyc_state_update_14_port, 
               Z(13) => cyc_state_update_13_port, Z(12) => 
               cyc_state_update_12_port, Z(11) => cyc_state_update_11_port, 
               Z(10) => cyc_state_update_10_port, Z(9) => 
               cyc_state_update_9_port, Z(8) => cyc_state_update_8_port, Z(7) 
               => cyc_state_update_7_port, Z(6) => cyc_state_update_6_port, 
               Z(5) => cyc_state_update_5_port, Z(4) => cyc_state_update_4_port
               , Z(3) => cyc_state_update_3_port, Z(2) => 
               cyc_state_update_2_port, Z(1) => cyc_state_update_1_port, Z(0) 
               => cyc_state_update_0_port );
   C1643_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 120 )
      port map(
         -- Connections to port 'DATA1'
         DATA(119) => state_main_out_plane2_127_port, DATA(118) => 
               state_main_out_plane2_126_port, DATA(117) => 
               state_main_out_plane2_125_port, DATA(116) => 
               state_main_out_plane2_124_port, DATA(115) => 
               state_main_out_plane2_123_port, DATA(114) => 
               state_main_out_plane2_122_port, DATA(113) => 
               state_main_out_plane2_121_port, DATA(112) => 
               state_main_out_plane2_120_port, DATA(111) => 
               state_main_out_plane2_119_port, DATA(110) => 
               state_main_out_plane2_118_port, DATA(109) => 
               state_main_out_plane2_117_port, DATA(108) => 
               state_main_out_plane2_116_port, DATA(107) => 
               state_main_out_plane2_115_port, DATA(106) => 
               state_main_out_plane2_114_port, DATA(105) => 
               state_main_out_plane2_113_port, DATA(104) => 
               state_main_out_plane2_112_port, DATA(103) => 
               state_main_out_plane2_111_port, DATA(102) => 
               state_main_out_plane2_110_port, DATA(101) => 
               state_main_out_plane2_109_port, DATA(100) => 
               state_main_out_plane2_108_port, DATA(99) => 
               state_main_out_plane2_107_port, DATA(98) => 
               state_main_out_plane2_106_port, DATA(97) => 
               state_main_out_plane2_105_port, DATA(96) => 
               state_main_out_plane2_104_port, DATA(95) => 
               state_main_out_plane2_103_port, DATA(94) => 
               state_main_out_plane2_102_port, DATA(93) => 
               state_main_out_plane2_101_port, DATA(92) => 
               state_main_out_plane2_100_port, DATA(91) => 
               state_main_out_plane2_99_port, DATA(90) => 
               state_main_out_plane2_98_port, DATA(89) => 
               state_main_out_plane2_97_port, DATA(88) => 
               state_main_out_plane2_96_port, DATA(87) => 
               state_main_out_plane2_95_port, DATA(86) => 
               state_main_out_plane2_94_port, DATA(85) => 
               state_main_out_plane2_93_port, DATA(84) => 
               state_main_out_plane2_92_port, DATA(83) => 
               state_main_out_plane2_91_port, DATA(82) => 
               state_main_out_plane2_90_port, DATA(81) => 
               state_main_out_plane2_89_port, DATA(80) => 
               state_main_out_plane2_88_port, DATA(79) => 
               state_main_out_plane2_87_port, DATA(78) => 
               state_main_out_plane2_86_port, DATA(77) => 
               state_main_out_plane2_85_port, DATA(76) => 
               state_main_out_plane2_84_port, DATA(75) => 
               state_main_out_plane2_83_port, DATA(74) => 
               state_main_out_plane2_82_port, DATA(73) => 
               state_main_out_plane2_81_port, DATA(72) => 
               state_main_out_plane2_80_port, DATA(71) => 
               state_main_out_plane2_79_port, DATA(70) => 
               state_main_out_plane2_78_port, DATA(69) => 
               state_main_out_plane2_77_port, DATA(68) => 
               state_main_out_plane2_76_port, DATA(67) => 
               state_main_out_plane2_75_port, DATA(66) => 
               state_main_out_plane2_74_port, DATA(65) => 
               state_main_out_plane2_73_port, DATA(64) => 
               state_main_out_plane2_72_port, DATA(63) => 
               state_main_out_plane2_71_port, DATA(62) => 
               state_main_out_plane2_70_port, DATA(61) => 
               state_main_out_plane2_69_port, DATA(60) => 
               state_main_out_plane2_68_port, DATA(59) => 
               state_main_out_plane2_67_port, DATA(58) => 
               state_main_out_plane2_66_port, DATA(57) => 
               state_main_out_plane2_65_port, DATA(56) => 
               state_main_out_plane2_64_port, DATA(55) => 
               state_main_out_plane2_63_port, DATA(54) => 
               state_main_out_plane2_62_port, DATA(53) => 
               state_main_out_plane2_61_port, DATA(52) => 
               state_main_out_plane2_60_port, DATA(51) => 
               state_main_out_plane2_59_port, DATA(50) => 
               state_main_out_plane2_58_port, DATA(49) => 
               state_main_out_plane2_57_port, DATA(48) => 
               state_main_out_plane2_56_port, DATA(47) => 
               state_main_out_plane2_55_port, DATA(46) => 
               state_main_out_plane2_54_port, DATA(45) => 
               state_main_out_plane2_53_port, DATA(44) => 
               state_main_out_plane2_52_port, DATA(43) => 
               state_main_out_plane2_51_port, DATA(42) => 
               state_main_out_plane2_50_port, DATA(41) => 
               state_main_out_plane2_49_port, DATA(40) => 
               state_main_out_plane2_48_port, DATA(39) => 
               state_main_out_plane2_47_port, DATA(38) => 
               state_main_out_plane2_46_port, DATA(37) => 
               state_main_out_plane2_45_port, DATA(36) => 
               state_main_out_plane2_44_port, DATA(35) => 
               state_main_out_plane2_43_port, DATA(34) => 
               state_main_out_plane2_42_port, DATA(33) => 
               state_main_out_plane2_41_port, DATA(32) => 
               state_main_out_plane2_40_port, DATA(31) => 
               state_main_out_plane2_39_port, DATA(30) => 
               state_main_out_plane2_38_port, DATA(29) => 
               state_main_out_plane2_37_port, DATA(28) => 
               state_main_out_plane2_36_port, DATA(27) => 
               state_main_out_plane2_35_port, DATA(26) => 
               state_main_out_plane2_34_port, DATA(25) => 
               state_main_out_plane2_33_port, DATA(24) => 
               state_main_out_plane2_32_port, DATA(23) => 
               state_main_out_plane2_23_port, DATA(22) => 
               state_main_out_plane2_22_port, DATA(21) => 
               state_main_out_plane2_21_port, DATA(20) => 
               state_main_out_plane2_20_port, DATA(19) => 
               state_main_out_plane2_19_port, DATA(18) => 
               state_main_out_plane2_18_port, DATA(17) => 
               state_main_out_plane2_17_port, DATA(16) => 
               state_main_out_plane2_16_port, DATA(15) => 
               state_main_out_plane2_15_port, DATA(14) => 
               state_main_out_plane2_14_port, DATA(13) => 
               state_main_out_plane2_13_port, DATA(12) => 
               state_main_out_plane2_12_port, DATA(11) => 
               state_main_out_plane2_11_port, DATA(10) => 
               state_main_out_plane2_10_port, DATA(9) => 
               state_main_out_plane2_9_port, DATA(8) => 
               state_main_out_plane2_8_port, DATA(7) => 
               state_main_out_plane2_7_port, DATA(6) => 
               state_main_out_plane2_6_port, DATA(5) => 
               state_main_out_plane2_5_port, DATA(4) => 
               state_main_out_plane2_4_port, DATA(3) => 
               state_main_out_plane2_3_port, DATA(2) => 
               state_main_out_plane2_2_port, DATA(1) => 
               state_main_out_plane2_1_port, DATA(0) => 
               state_main_out_plane2_0_port, 
         -- Connections to port 'DATA2'
         DATA(239) => cyc_state_update_127_port, DATA(238) => 
               cyc_state_update_126_port, DATA(237) => 
               cyc_state_update_125_port, DATA(236) => 
               cyc_state_update_124_port, DATA(235) => 
               cyc_state_update_123_port, DATA(234) => 
               cyc_state_update_122_port, DATA(233) => 
               cyc_state_update_121_port, DATA(232) => 
               cyc_state_update_120_port, DATA(231) => 
               cyc_state_update_119_port, DATA(230) => 
               cyc_state_update_118_port, DATA(229) => 
               cyc_state_update_117_port, DATA(228) => 
               cyc_state_update_116_port, DATA(227) => 
               cyc_state_update_115_port, DATA(226) => 
               cyc_state_update_114_port, DATA(225) => 
               cyc_state_update_113_port, DATA(224) => 
               cyc_state_update_112_port, DATA(223) => 
               cyc_state_update_111_port, DATA(222) => 
               cyc_state_update_110_port, DATA(221) => 
               cyc_state_update_109_port, DATA(220) => 
               cyc_state_update_108_port, DATA(219) => 
               cyc_state_update_107_port, DATA(218) => 
               cyc_state_update_106_port, DATA(217) => 
               cyc_state_update_105_port, DATA(216) => 
               cyc_state_update_104_port, DATA(215) => 
               cyc_state_update_103_port, DATA(214) => 
               cyc_state_update_102_port, DATA(213) => 
               cyc_state_update_101_port, DATA(212) => 
               cyc_state_update_100_port, DATA(211) => cyc_state_update_99_port
               , DATA(210) => cyc_state_update_98_port, DATA(209) => 
               cyc_state_update_97_port, DATA(208) => cyc_state_update_96_port,
               DATA(207) => cyc_state_update_95_port, DATA(206) => 
               cyc_state_update_94_port, DATA(205) => cyc_state_update_93_port,
               DATA(204) => cyc_state_update_92_port, DATA(203) => 
               cyc_state_update_91_port, DATA(202) => cyc_state_update_90_port,
               DATA(201) => cyc_state_update_89_port, DATA(200) => 
               cyc_state_update_88_port, DATA(199) => cyc_state_update_87_port,
               DATA(198) => cyc_state_update_86_port, DATA(197) => 
               cyc_state_update_85_port, DATA(196) => cyc_state_update_84_port,
               DATA(195) => cyc_state_update_83_port, DATA(194) => 
               cyc_state_update_82_port, DATA(193) => cyc_state_update_81_port,
               DATA(192) => cyc_state_update_80_port, DATA(191) => 
               cyc_state_update_79_port, DATA(190) => cyc_state_update_78_port,
               DATA(189) => cyc_state_update_77_port, DATA(188) => 
               cyc_state_update_76_port, DATA(187) => cyc_state_update_75_port,
               DATA(186) => cyc_state_update_74_port, DATA(185) => 
               cyc_state_update_73_port, DATA(184) => cyc_state_update_72_port,
               DATA(183) => cyc_state_update_71_port, DATA(182) => 
               cyc_state_update_70_port, DATA(181) => cyc_state_update_69_port,
               DATA(180) => cyc_state_update_68_port, DATA(179) => 
               cyc_state_update_67_port, DATA(178) => cyc_state_update_66_port,
               DATA(177) => cyc_state_update_65_port, DATA(176) => 
               cyc_state_update_64_port, DATA(175) => cyc_state_update_63_port,
               DATA(174) => cyc_state_update_62_port, DATA(173) => 
               cyc_state_update_61_port, DATA(172) => cyc_state_update_60_port,
               DATA(171) => cyc_state_update_59_port, DATA(170) => 
               cyc_state_update_58_port, DATA(169) => cyc_state_update_57_port,
               DATA(168) => cyc_state_update_56_port, DATA(167) => 
               cyc_state_update_55_port, DATA(166) => cyc_state_update_54_port,
               DATA(165) => cyc_state_update_53_port, DATA(164) => 
               cyc_state_update_52_port, DATA(163) => cyc_state_update_51_port,
               DATA(162) => cyc_state_update_50_port, DATA(161) => 
               cyc_state_update_49_port, DATA(160) => cyc_state_update_48_port,
               DATA(159) => cyc_state_update_47_port, DATA(158) => 
               cyc_state_update_46_port, DATA(157) => cyc_state_update_45_port,
               DATA(156) => cyc_state_update_44_port, DATA(155) => 
               cyc_state_update_43_port, DATA(154) => cyc_state_update_42_port,
               DATA(153) => cyc_state_update_41_port, DATA(152) => 
               cyc_state_update_40_port, DATA(151) => cyc_state_update_39_port,
               DATA(150) => cyc_state_update_38_port, DATA(149) => 
               cyc_state_update_37_port, DATA(148) => cyc_state_update_36_port,
               DATA(147) => cyc_state_update_35_port, DATA(146) => 
               cyc_state_update_34_port, DATA(145) => cyc_state_update_33_port,
               DATA(144) => cyc_state_update_32_port, DATA(143) => 
               cyc_state_update_23_port, DATA(142) => cyc_state_update_22_port,
               DATA(141) => cyc_state_update_21_port, DATA(140) => 
               cyc_state_update_20_port, DATA(139) => cyc_state_update_19_port,
               DATA(138) => cyc_state_update_18_port, DATA(137) => 
               cyc_state_update_17_port, DATA(136) => cyc_state_update_16_port,
               DATA(135) => cyc_state_update_15_port, DATA(134) => 
               cyc_state_update_14_port, DATA(133) => cyc_state_update_13_port,
               DATA(132) => cyc_state_update_12_port, DATA(131) => 
               cyc_state_update_11_port, DATA(130) => cyc_state_update_10_port,
               DATA(129) => cyc_state_update_9_port, DATA(128) => 
               cyc_state_update_8_port, DATA(127) => cyc_state_update_7_port, 
               DATA(126) => cyc_state_update_6_port, DATA(125) => 
               cyc_state_update_5_port, DATA(124) => cyc_state_update_4_port, 
               DATA(123) => cyc_state_update_3_port, DATA(122) => 
               cyc_state_update_2_port, DATA(121) => cyc_state_update_1_port, 
               DATA(120) => cyc_state_update_0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N18, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N19, 
         -- Connections to port 'Z'
         Z(119) => plane_2_input_127_port, Z(118) => plane_2_input_126_port, 
               Z(117) => plane_2_input_125_port, Z(116) => 
               plane_2_input_124_port, Z(115) => plane_2_input_123_port, Z(114)
               => plane_2_input_122_port, Z(113) => plane_2_input_121_port, 
               Z(112) => plane_2_input_120_port, Z(111) => 
               plane_2_input_119_port, Z(110) => plane_2_input_118_port, Z(109)
               => plane_2_input_117_port, Z(108) => plane_2_input_116_port, 
               Z(107) => plane_2_input_115_port, Z(106) => 
               plane_2_input_114_port, Z(105) => plane_2_input_113_port, Z(104)
               => plane_2_input_112_port, Z(103) => plane_2_input_111_port, 
               Z(102) => plane_2_input_110_port, Z(101) => 
               plane_2_input_109_port, Z(100) => plane_2_input_108_port, Z(99) 
               => plane_2_input_107_port, Z(98) => plane_2_input_106_port, 
               Z(97) => plane_2_input_105_port, Z(96) => plane_2_input_104_port
               , Z(95) => plane_2_input_103_port, Z(94) => 
               plane_2_input_102_port, Z(93) => plane_2_input_101_port, Z(92) 
               => plane_2_input_100_port, Z(91) => plane_2_input_99_port, Z(90)
               => plane_2_input_98_port, Z(89) => plane_2_input_97_port, Z(88) 
               => plane_2_input_96_port, Z(87) => plane_2_input_95_port, Z(86) 
               => plane_2_input_94_port, Z(85) => plane_2_input_93_port, Z(84) 
               => plane_2_input_92_port, Z(83) => plane_2_input_91_port, Z(82) 
               => plane_2_input_90_port, Z(81) => plane_2_input_89_port, Z(80) 
               => plane_2_input_88_port, Z(79) => plane_2_input_87_port, Z(78) 
               => plane_2_input_86_port, Z(77) => plane_2_input_85_port, Z(76) 
               => plane_2_input_84_port, Z(75) => plane_2_input_83_port, Z(74) 
               => plane_2_input_82_port, Z(73) => plane_2_input_81_port, Z(72) 
               => plane_2_input_80_port, Z(71) => plane_2_input_79_port, Z(70) 
               => plane_2_input_78_port, Z(69) => plane_2_input_77_port, Z(68) 
               => plane_2_input_76_port, Z(67) => plane_2_input_75_port, Z(66) 
               => plane_2_input_74_port, Z(65) => plane_2_input_73_port, Z(64) 
               => plane_2_input_72_port, Z(63) => plane_2_input_71_port, Z(62) 
               => plane_2_input_70_port, Z(61) => plane_2_input_69_port, Z(60) 
               => plane_2_input_68_port, Z(59) => plane_2_input_67_port, Z(58) 
               => plane_2_input_66_port, Z(57) => plane_2_input_65_port, Z(56) 
               => plane_2_input_64_port, Z(55) => plane_2_input_63_port, Z(54) 
               => plane_2_input_62_port, Z(53) => plane_2_input_61_port, Z(52) 
               => plane_2_input_60_port, Z(51) => plane_2_input_59_port, Z(50) 
               => plane_2_input_58_port, Z(49) => plane_2_input_57_port, Z(48) 
               => plane_2_input_56_port, Z(47) => plane_2_input_55_port, Z(46) 
               => plane_2_input_54_port, Z(45) => plane_2_input_53_port, Z(44) 
               => plane_2_input_52_port, Z(43) => plane_2_input_51_port, Z(42) 
               => plane_2_input_50_port, Z(41) => plane_2_input_49_port, Z(40) 
               => plane_2_input_48_port, Z(39) => plane_2_input_47_port, Z(38) 
               => plane_2_input_46_port, Z(37) => plane_2_input_45_port, Z(36) 
               => plane_2_input_44_port, Z(35) => plane_2_input_43_port, Z(34) 
               => plane_2_input_42_port, Z(33) => plane_2_input_41_port, Z(32) 
               => plane_2_input_40_port, Z(31) => plane_2_input_39_port, Z(30) 
               => plane_2_input_38_port, Z(29) => plane_2_input_37_port, Z(28) 
               => plane_2_input_36_port, Z(27) => plane_2_input_35_port, Z(26) 
               => plane_2_input_34_port, Z(25) => plane_2_input_33_port, Z(24) 
               => plane_2_input_32_port, Z(23) => plane_2_input_23, Z(22) => 
               plane_2_input_22, Z(21) => plane_2_input_21, Z(20) => 
               plane_2_input_20, Z(19) => plane_2_input_19, Z(18) => 
               plane_2_input_18, Z(17) => plane_2_input_17, Z(16) => 
               plane_2_input_16, Z(15) => plane_2_input_15, Z(14) => 
               plane_2_input_14, Z(13) => plane_2_input_13, Z(12) => 
               plane_2_input_12, Z(11) => plane_2_input_11, Z(10) => 
               plane_2_input_10, Z(9) => plane_2_input_9, Z(8) => 
               plane_2_input_8, Z(7) => plane_2_input_7, Z(6) => 
               plane_2_input_6, Z(5) => plane_2_input_5, Z(4) => 
               plane_2_input_4, Z(3) => plane_2_input_3, Z(2) => 
               plane_2_input_2, Z(1) => plane_2_input_1, Z(0) => 
               plane_2_input_0 );
   B_18 : GTECH_BUF port map( A => N574, Z => N18);
   B_19 : GTECH_BUF port map( A => state_main_sel(6), Z => N19);
   C1644_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 128 )
      port map(
         -- Connections to port 'DATA1'
         DATA(127) => cyc_state_update_127_port, DATA(126) => 
               cyc_state_update_126_port, DATA(125) => 
               cyc_state_update_125_port, DATA(124) => 
               cyc_state_update_124_port, DATA(123) => 
               cyc_state_update_123_port, DATA(122) => 
               cyc_state_update_122_port, DATA(121) => 
               cyc_state_update_121_port, DATA(120) => 
               cyc_state_update_120_port, DATA(119) => 
               cyc_state_update_119_port, DATA(118) => 
               cyc_state_update_118_port, DATA(117) => 
               cyc_state_update_117_port, DATA(116) => 
               cyc_state_update_116_port, DATA(115) => 
               cyc_state_update_115_port, DATA(114) => 
               cyc_state_update_114_port, DATA(113) => 
               cyc_state_update_113_port, DATA(112) => 
               cyc_state_update_112_port, DATA(111) => 
               cyc_state_update_111_port, DATA(110) => 
               cyc_state_update_110_port, DATA(109) => 
               cyc_state_update_109_port, DATA(108) => 
               cyc_state_update_108_port, DATA(107) => 
               cyc_state_update_107_port, DATA(106) => 
               cyc_state_update_106_port, DATA(105) => 
               cyc_state_update_105_port, DATA(104) => 
               cyc_state_update_104_port, DATA(103) => 
               cyc_state_update_103_port, DATA(102) => 
               cyc_state_update_102_port, DATA(101) => 
               cyc_state_update_101_port, DATA(100) => 
               cyc_state_update_100_port, DATA(99) => cyc_state_update_99_port,
               DATA(98) => cyc_state_update_98_port, DATA(97) => 
               cyc_state_update_97_port, DATA(96) => cyc_state_update_96_port, 
               DATA(95) => cyc_state_update_95_port, DATA(94) => 
               cyc_state_update_94_port, DATA(93) => cyc_state_update_93_port, 
               DATA(92) => cyc_state_update_92_port, DATA(91) => 
               cyc_state_update_91_port, DATA(90) => cyc_state_update_90_port, 
               DATA(89) => cyc_state_update_89_port, DATA(88) => 
               cyc_state_update_88_port, DATA(87) => cyc_state_update_87_port, 
               DATA(86) => cyc_state_update_86_port, DATA(85) => 
               cyc_state_update_85_port, DATA(84) => cyc_state_update_84_port, 
               DATA(83) => cyc_state_update_83_port, DATA(82) => 
               cyc_state_update_82_port, DATA(81) => cyc_state_update_81_port, 
               DATA(80) => cyc_state_update_80_port, DATA(79) => 
               cyc_state_update_79_port, DATA(78) => cyc_state_update_78_port, 
               DATA(77) => cyc_state_update_77_port, DATA(76) => 
               cyc_state_update_76_port, DATA(75) => cyc_state_update_75_port, 
               DATA(74) => cyc_state_update_74_port, DATA(73) => 
               cyc_state_update_73_port, DATA(72) => cyc_state_update_72_port, 
               DATA(71) => cyc_state_update_71_port, DATA(70) => 
               cyc_state_update_70_port, DATA(69) => cyc_state_update_69_port, 
               DATA(68) => cyc_state_update_68_port, DATA(67) => 
               cyc_state_update_67_port, DATA(66) => cyc_state_update_66_port, 
               DATA(65) => cyc_state_update_65_port, DATA(64) => 
               cyc_state_update_64_port, DATA(63) => cyc_state_update_63_port, 
               DATA(62) => cyc_state_update_62_port, DATA(61) => 
               cyc_state_update_61_port, DATA(60) => cyc_state_update_60_port, 
               DATA(59) => cyc_state_update_59_port, DATA(58) => 
               cyc_state_update_58_port, DATA(57) => cyc_state_update_57_port, 
               DATA(56) => cyc_state_update_56_port, DATA(55) => 
               cyc_state_update_55_port, DATA(54) => cyc_state_update_54_port, 
               DATA(53) => cyc_state_update_53_port, DATA(52) => 
               cyc_state_update_52_port, DATA(51) => cyc_state_update_51_port, 
               DATA(50) => cyc_state_update_50_port, DATA(49) => 
               cyc_state_update_49_port, DATA(48) => cyc_state_update_48_port, 
               DATA(47) => cyc_state_update_47_port, DATA(46) => 
               cyc_state_update_46_port, DATA(45) => cyc_state_update_45_port, 
               DATA(44) => cyc_state_update_44_port, DATA(43) => 
               cyc_state_update_43_port, DATA(42) => cyc_state_update_42_port, 
               DATA(41) => cyc_state_update_41_port, DATA(40) => 
               cyc_state_update_40_port, DATA(39) => cyc_state_update_39_port, 
               DATA(38) => cyc_state_update_38_port, DATA(37) => 
               cyc_state_update_37_port, DATA(36) => cyc_state_update_36_port, 
               DATA(35) => cyc_state_update_35_port, DATA(34) => 
               cyc_state_update_34_port, DATA(33) => cyc_state_update_33_port, 
               DATA(32) => cyc_state_update_32_port, DATA(31) => 
               cyc_state_update_31_port, DATA(30) => cyc_state_update_30_port, 
               DATA(29) => cyc_state_update_29_port, DATA(28) => 
               cyc_state_update_28_port, DATA(27) => cyc_state_update_27_port, 
               DATA(26) => cyc_state_update_26_port, DATA(25) => 
               cyc_state_update_25_port, DATA(24) => cyc_state_update_24_port, 
               DATA(23) => cyc_state_update_23_port, DATA(22) => 
               cyc_state_update_22_port, DATA(21) => cyc_state_update_21_port, 
               DATA(20) => cyc_state_update_20_port, DATA(19) => 
               cyc_state_update_19_port, DATA(18) => cyc_state_update_18_port, 
               DATA(17) => cyc_state_update_17_port, DATA(16) => 
               cyc_state_update_16_port, DATA(15) => cyc_state_update_15_port, 
               DATA(14) => cyc_state_update_14_port, DATA(13) => 
               cyc_state_update_13_port, DATA(12) => cyc_state_update_12_port, 
               DATA(11) => cyc_state_update_11_port, DATA(10) => 
               cyc_state_update_10_port, DATA(9) => cyc_state_update_9_port, 
               DATA(8) => cyc_state_update_8_port, DATA(7) => 
               cyc_state_update_7_port, DATA(6) => cyc_state_update_6_port, 
               DATA(5) => cyc_state_update_5_port, DATA(4) => 
               cyc_state_update_4_port, DATA(3) => cyc_state_update_3_port, 
               DATA(2) => cyc_state_update_2_port, DATA(1) => 
               cyc_state_update_1_port, DATA(0) => cyc_state_update_0_port, 
         -- Connections to port 'DATA2'
         DATA(255) => perm_output_127_port, DATA(254) => perm_output_126_port, 
               DATA(253) => perm_output_125_port, DATA(252) => 
               perm_output_124_port, DATA(251) => perm_output_123_port, 
               DATA(250) => perm_output_122_port, DATA(249) => 
               perm_output_121_port, DATA(248) => perm_output_120_port, 
               DATA(247) => perm_output_119_port, DATA(246) => 
               perm_output_118_port, DATA(245) => perm_output_117_port, 
               DATA(244) => perm_output_116_port, DATA(243) => 
               perm_output_115_port, DATA(242) => perm_output_114_port, 
               DATA(241) => perm_output_113_port, DATA(240) => 
               perm_output_112_port, DATA(239) => perm_output_111_port, 
               DATA(238) => perm_output_110_port, DATA(237) => 
               perm_output_109_port, DATA(236) => perm_output_108_port, 
               DATA(235) => perm_output_107_port, DATA(234) => 
               perm_output_106_port, DATA(233) => perm_output_105_port, 
               DATA(232) => perm_output_104_port, DATA(231) => 
               perm_output_103_port, DATA(230) => perm_output_102_port, 
               DATA(229) => perm_output_101_port, DATA(228) => 
               perm_output_100_port, DATA(227) => perm_output_99_port, 
               DATA(226) => perm_output_98_port, DATA(225) => 
               perm_output_97_port, DATA(224) => perm_output_96_port, DATA(223)
               => perm_output_95_port, DATA(222) => perm_output_94_port, 
               DATA(221) => perm_output_93_port, DATA(220) => 
               perm_output_92_port, DATA(219) => perm_output_91_port, DATA(218)
               => perm_output_90_port, DATA(217) => perm_output_89_port, 
               DATA(216) => perm_output_88_port, DATA(215) => 
               perm_output_87_port, DATA(214) => perm_output_86_port, DATA(213)
               => perm_output_85_port, DATA(212) => perm_output_84_port, 
               DATA(211) => perm_output_83_port, DATA(210) => 
               perm_output_82_port, DATA(209) => perm_output_81_port, DATA(208)
               => perm_output_80_port, DATA(207) => perm_output_79_port, 
               DATA(206) => perm_output_78_port, DATA(205) => 
               perm_output_77_port, DATA(204) => perm_output_76_port, DATA(203)
               => perm_output_75_port, DATA(202) => perm_output_74_port, 
               DATA(201) => perm_output_73_port, DATA(200) => 
               perm_output_72_port, DATA(199) => perm_output_71_port, DATA(198)
               => perm_output_70_port, DATA(197) => perm_output_69_port, 
               DATA(196) => perm_output_68_port, DATA(195) => 
               perm_output_67_port, DATA(194) => perm_output_66_port, DATA(193)
               => perm_output_65_port, DATA(192) => perm_output_64_port, 
               DATA(191) => perm_output_63_port, DATA(190) => 
               perm_output_62_port, DATA(189) => perm_output_61_port, DATA(188)
               => perm_output_60_port, DATA(187) => perm_output_59_port, 
               DATA(186) => perm_output_58_port, DATA(185) => 
               perm_output_57_port, DATA(184) => perm_output_56_port, DATA(183)
               => perm_output_55_port, DATA(182) => perm_output_54_port, 
               DATA(181) => perm_output_53_port, DATA(180) => 
               perm_output_52_port, DATA(179) => perm_output_51_port, DATA(178)
               => perm_output_50_port, DATA(177) => perm_output_49_port, 
               DATA(176) => perm_output_48_port, DATA(175) => 
               perm_output_47_port, DATA(174) => perm_output_46_port, DATA(173)
               => perm_output_45_port, DATA(172) => perm_output_44_port, 
               DATA(171) => perm_output_43_port, DATA(170) => 
               perm_output_42_port, DATA(169) => perm_output_41_port, DATA(168)
               => perm_output_40_port, DATA(167) => perm_output_39_port, 
               DATA(166) => perm_output_38_port, DATA(165) => 
               perm_output_37_port, DATA(164) => perm_output_36_port, DATA(163)
               => perm_output_35_port, DATA(162) => perm_output_34_port, 
               DATA(161) => perm_output_33_port, DATA(160) => 
               perm_output_32_port, DATA(159) => perm_output_31_port, DATA(158)
               => perm_output_30_port, DATA(157) => perm_output_29_port, 
               DATA(156) => perm_output_28_port, DATA(155) => 
               perm_output_27_port, DATA(154) => perm_output_26_port, DATA(153)
               => perm_output_25_port, DATA(152) => perm_output_24_port, 
               DATA(151) => perm_output_23_port, DATA(150) => 
               perm_output_22_port, DATA(149) => perm_output_21_port, DATA(148)
               => perm_output_20_port, DATA(147) => perm_output_19_port, 
               DATA(146) => perm_output_18_port, DATA(145) => 
               perm_output_17_port, DATA(144) => perm_output_16_port, DATA(143)
               => perm_output_15_port, DATA(142) => perm_output_14_port, 
               DATA(141) => perm_output_13_port, DATA(140) => 
               perm_output_12_port, DATA(139) => perm_output_11_port, DATA(138)
               => perm_output_10_port, DATA(137) => perm_output_9_port, 
               DATA(136) => perm_output_8_port, DATA(135) => perm_output_7_port
               , DATA(134) => perm_output_6_port, DATA(133) => 
               perm_output_5_port, DATA(132) => perm_output_4_port, DATA(131) 
               => perm_output_3_port, DATA(130) => perm_output_2_port, 
               DATA(129) => perm_output_1_port, DATA(128) => perm_output_0_port
               , 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N20, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N21, 
         -- Connections to port 'Z'
         Z(127) => N310, Z(126) => N309, Z(125) => N308, Z(124) => N307, Z(123)
               => N306, Z(122) => N305, Z(121) => N304, Z(120) => N303, Z(119) 
               => N302, Z(118) => N301, Z(117) => N300, Z(116) => N299, Z(115) 
               => N298, Z(114) => N297, Z(113) => N296, Z(112) => N295, Z(111) 
               => N294, Z(110) => N293, Z(109) => N292, Z(108) => N291, Z(107) 
               => N290, Z(106) => N289, Z(105) => N288, Z(104) => N287, Z(103) 
               => N286, Z(102) => N285, Z(101) => N284, Z(100) => N283, Z(99) 
               => N282, Z(98) => N281, Z(97) => N280, Z(96) => N279, Z(95) => 
               N278, Z(94) => N277, Z(93) => N276, Z(92) => N275, Z(91) => N274
               , Z(90) => N273, Z(89) => N272, Z(88) => N271, Z(87) => N270, 
               Z(86) => N269, Z(85) => N268, Z(84) => N267, Z(83) => N266, 
               Z(82) => N265, Z(81) => N264, Z(80) => N263, Z(79) => N262, 
               Z(78) => N261, Z(77) => N260, Z(76) => N259, Z(75) => N258, 
               Z(74) => N257, Z(73) => N256, Z(72) => N255, Z(71) => N254, 
               Z(70) => N253, Z(69) => N252, Z(68) => N251, Z(67) => N250, 
               Z(66) => N249, Z(65) => N248, Z(64) => N247, Z(63) => N246, 
               Z(62) => N245, Z(61) => N244, Z(60) => N243, Z(59) => N242, 
               Z(58) => N241, Z(57) => N240, Z(56) => N239, Z(55) => N238, 
               Z(54) => N237, Z(53) => N236, Z(52) => N235, Z(51) => N234, 
               Z(50) => N233, Z(49) => N232, Z(48) => N231, Z(47) => N230, 
               Z(46) => N229, Z(45) => N228, Z(44) => N227, Z(43) => N226, 
               Z(42) => N225, Z(41) => N224, Z(40) => N223, Z(39) => N222, 
               Z(38) => N221, Z(37) => N220, Z(36) => N219, Z(35) => N218, 
               Z(34) => N217, Z(33) => N216, Z(32) => N215, Z(31) => N214, 
               Z(30) => N213, Z(29) => N212, Z(28) => N211, Z(27) => N210, 
               Z(26) => N209, Z(25) => N208, Z(24) => N207, Z(23) => N206, 
               Z(22) => N205, Z(21) => N204, Z(20) => N203, Z(19) => N202, 
               Z(18) => N201, Z(17) => N200, Z(16) => N199, Z(15) => N198, 
               Z(14) => N197, Z(13) => N196, Z(12) => N195, Z(11) => N194, 
               Z(10) => N193, Z(9) => N192, Z(8) => N191, Z(7) => N190, Z(6) =>
               N189, Z(5) => N188, Z(4) => N187, Z(3) => N186, Z(2) => N185, 
               Z(1) => N184, Z(0) => N183 );
   B_20 : GTECH_BUF port map( A => N182, Z => N20);
   B_21 : GTECH_BUF port map( A => state_main_sel(0), Z => N21);
   C1645_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 128 )
      port map(
         -- Connections to port 'DATA1'
         DATA(127) => N310, DATA(126) => N309, DATA(125) => N308, DATA(124) => 
               N307, DATA(123) => N306, DATA(122) => N305, DATA(121) => N304, 
               DATA(120) => N303, DATA(119) => N302, DATA(118) => N301, 
               DATA(117) => N300, DATA(116) => N299, DATA(115) => N298, 
               DATA(114) => N297, DATA(113) => N296, DATA(112) => N295, 
               DATA(111) => N294, DATA(110) => N293, DATA(109) => N292, 
               DATA(108) => N291, DATA(107) => N290, DATA(106) => N289, 
               DATA(105) => N288, DATA(104) => N287, DATA(103) => N286, 
               DATA(102) => N285, DATA(101) => N284, DATA(100) => N283, 
               DATA(99) => N282, DATA(98) => N281, DATA(97) => N280, DATA(96) 
               => N279, DATA(95) => N278, DATA(94) => N277, DATA(93) => N276, 
               DATA(92) => N275, DATA(91) => N274, DATA(90) => N273, DATA(89) 
               => N272, DATA(88) => N271, DATA(87) => N270, DATA(86) => N269, 
               DATA(85) => N268, DATA(84) => N267, DATA(83) => N266, DATA(82) 
               => N265, DATA(81) => N264, DATA(80) => N263, DATA(79) => N262, 
               DATA(78) => N261, DATA(77) => N260, DATA(76) => N259, DATA(75) 
               => N258, DATA(74) => N257, DATA(73) => N256, DATA(72) => N255, 
               DATA(71) => N254, DATA(70) => N253, DATA(69) => N252, DATA(68) 
               => N251, DATA(67) => N250, DATA(66) => N249, DATA(65) => N248, 
               DATA(64) => N247, DATA(63) => N246, DATA(62) => N245, DATA(61) 
               => N244, DATA(60) => N243, DATA(59) => N242, DATA(58) => N241, 
               DATA(57) => N240, DATA(56) => N239, DATA(55) => N238, DATA(54) 
               => N237, DATA(53) => N236, DATA(52) => N235, DATA(51) => N234, 
               DATA(50) => N233, DATA(49) => N232, DATA(48) => N231, DATA(47) 
               => N230, DATA(46) => N229, DATA(45) => N228, DATA(44) => N227, 
               DATA(43) => N226, DATA(42) => N225, DATA(41) => N224, DATA(40) 
               => N223, DATA(39) => N222, DATA(38) => N221, DATA(37) => N220, 
               DATA(36) => N219, DATA(35) => N218, DATA(34) => N217, DATA(33) 
               => N216, DATA(32) => N215, DATA(31) => N214, DATA(30) => N213, 
               DATA(29) => N212, DATA(28) => N211, DATA(27) => N210, DATA(26) 
               => N209, DATA(25) => N208, DATA(24) => N207, DATA(23) => N206, 
               DATA(22) => N205, DATA(21) => N204, DATA(20) => N203, DATA(19) 
               => N202, DATA(18) => N201, DATA(17) => N200, DATA(16) => N199, 
               DATA(15) => N198, DATA(14) => N197, DATA(13) => N196, DATA(12) 
               => N195, DATA(11) => N194, DATA(10) => N193, DATA(9) => N192, 
               DATA(8) => N191, DATA(7) => N190, DATA(6) => N189, DATA(5) => 
               N188, DATA(4) => N187, DATA(3) => N186, DATA(2) => N185, DATA(1)
               => N184, DATA(0) => N183, 
         -- Connections to port 'DATA2'
         DATA(255) => X_Logic0_port, DATA(254) => X_Logic0_port, DATA(253) => 
               X_Logic0_port, DATA(252) => X_Logic0_port, DATA(251) => 
               X_Logic0_port, DATA(250) => X_Logic0_port, DATA(249) => 
               X_Logic0_port, DATA(248) => X_Logic0_port, DATA(247) => 
               X_Logic0_port, DATA(246) => X_Logic0_port, DATA(245) => 
               X_Logic0_port, DATA(244) => X_Logic0_port, DATA(243) => 
               X_Logic0_port, DATA(242) => X_Logic0_port, DATA(241) => 
               X_Logic0_port, DATA(240) => X_Logic0_port, DATA(239) => 
               X_Logic0_port, DATA(238) => X_Logic0_port, DATA(237) => 
               X_Logic0_port, DATA(236) => X_Logic0_port, DATA(235) => 
               X_Logic0_port, DATA(234) => X_Logic0_port, DATA(233) => 
               X_Logic0_port, DATA(232) => X_Logic0_port, DATA(231) => 
               X_Logic0_port, DATA(230) => X_Logic0_port, DATA(229) => 
               X_Logic0_port, DATA(228) => X_Logic0_port, DATA(227) => 
               X_Logic0_port, DATA(226) => X_Logic0_port, DATA(225) => 
               X_Logic0_port, DATA(224) => X_Logic0_port, DATA(223) => 
               X_Logic0_port, DATA(222) => X_Logic0_port, DATA(221) => 
               X_Logic0_port, DATA(220) => X_Logic0_port, DATA(219) => 
               X_Logic0_port, DATA(218) => X_Logic0_port, DATA(217) => 
               X_Logic0_port, DATA(216) => X_Logic0_port, DATA(215) => 
               X_Logic0_port, DATA(214) => X_Logic0_port, DATA(213) => 
               X_Logic0_port, DATA(212) => X_Logic0_port, DATA(211) => 
               X_Logic0_port, DATA(210) => X_Logic0_port, DATA(209) => 
               X_Logic0_port, DATA(208) => X_Logic0_port, DATA(207) => 
               X_Logic0_port, DATA(206) => X_Logic0_port, DATA(205) => 
               X_Logic0_port, DATA(204) => X_Logic0_port, DATA(203) => 
               X_Logic0_port, DATA(202) => X_Logic0_port, DATA(201) => 
               X_Logic0_port, DATA(200) => X_Logic0_port, DATA(199) => 
               X_Logic0_port, DATA(198) => X_Logic0_port, DATA(197) => 
               X_Logic0_port, DATA(196) => X_Logic0_port, DATA(195) => 
               X_Logic0_port, DATA(194) => X_Logic0_port, DATA(193) => 
               X_Logic0_port, DATA(192) => X_Logic0_port, DATA(191) => 
               X_Logic0_port, DATA(190) => X_Logic0_port, DATA(189) => 
               X_Logic0_port, DATA(188) => X_Logic0_port, DATA(187) => 
               X_Logic0_port, DATA(186) => X_Logic0_port, DATA(185) => 
               X_Logic0_port, DATA(184) => X_Logic0_port, DATA(183) => 
               X_Logic0_port, DATA(182) => X_Logic0_port, DATA(181) => 
               X_Logic0_port, DATA(180) => X_Logic0_port, DATA(179) => 
               X_Logic0_port, DATA(178) => X_Logic0_port, DATA(177) => 
               X_Logic0_port, DATA(176) => X_Logic0_port, DATA(175) => 
               X_Logic0_port, DATA(174) => X_Logic0_port, DATA(173) => 
               X_Logic0_port, DATA(172) => X_Logic0_port, DATA(171) => 
               X_Logic0_port, DATA(170) => X_Logic0_port, DATA(169) => 
               X_Logic0_port, DATA(168) => X_Logic0_port, DATA(167) => 
               X_Logic0_port, DATA(166) => X_Logic0_port, DATA(165) => 
               X_Logic0_port, DATA(164) => X_Logic0_port, DATA(163) => 
               X_Logic0_port, DATA(162) => X_Logic0_port, DATA(161) => 
               X_Logic0_port, DATA(160) => X_Logic0_port, DATA(159) => 
               X_Logic0_port, DATA(158) => X_Logic0_port, DATA(157) => 
               X_Logic0_port, DATA(156) => X_Logic0_port, DATA(155) => 
               X_Logic0_port, DATA(154) => X_Logic0_port, DATA(153) => 
               X_Logic0_port, DATA(152) => X_Logic0_port, DATA(151) => 
               X_Logic0_port, DATA(150) => X_Logic0_port, DATA(149) => 
               X_Logic0_port, DATA(148) => X_Logic0_port, DATA(147) => 
               X_Logic0_port, DATA(146) => X_Logic0_port, DATA(145) => 
               X_Logic0_port, DATA(144) => X_Logic0_port, DATA(143) => 
               X_Logic0_port, DATA(142) => X_Logic0_port, DATA(141) => 
               X_Logic0_port, DATA(140) => X_Logic0_port, DATA(139) => 
               X_Logic0_port, DATA(138) => X_Logic0_port, DATA(137) => 
               X_Logic0_port, DATA(136) => X_Logic0_port, DATA(135) => 
               X_Logic0_port, DATA(134) => X_Logic0_port, DATA(133) => 
               X_Logic0_port, DATA(132) => X_Logic0_port, DATA(131) => 
               X_Logic0_port, DATA(130) => X_Logic0_port, DATA(129) => 
               X_Logic0_port, DATA(128) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N22, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N23, 
         -- Connections to port 'Z'
         Z(127) => state_main_in_p0_127_port, Z(126) => 
               state_main_in_p0_126_port, Z(125) => state_main_in_p0_125_port, 
               Z(124) => state_main_in_p0_124_port, Z(123) => 
               state_main_in_p0_123_port, Z(122) => state_main_in_p0_122_port, 
               Z(121) => state_main_in_p0_121_port, Z(120) => 
               state_main_in_p0_120_port, Z(119) => state_main_in_p0_119_port, 
               Z(118) => state_main_in_p0_118_port, Z(117) => 
               state_main_in_p0_117_port, Z(116) => state_main_in_p0_116_port, 
               Z(115) => state_main_in_p0_115_port, Z(114) => 
               state_main_in_p0_114_port, Z(113) => state_main_in_p0_113_port, 
               Z(112) => state_main_in_p0_112_port, Z(111) => 
               state_main_in_p0_111_port, Z(110) => state_main_in_p0_110_port, 
               Z(109) => state_main_in_p0_109_port, Z(108) => 
               state_main_in_p0_108_port, Z(107) => state_main_in_p0_107_port, 
               Z(106) => state_main_in_p0_106_port, Z(105) => 
               state_main_in_p0_105_port, Z(104) => state_main_in_p0_104_port, 
               Z(103) => state_main_in_p0_103_port, Z(102) => 
               state_main_in_p0_102_port, Z(101) => state_main_in_p0_101_port, 
               Z(100) => state_main_in_p0_100_port, Z(99) => 
               state_main_in_p0_99_port, Z(98) => state_main_in_p0_98_port, 
               Z(97) => state_main_in_p0_97_port, Z(96) => 
               state_main_in_p0_96_port, Z(95) => state_main_in_p0_95_port, 
               Z(94) => state_main_in_p0_94_port, Z(93) => 
               state_main_in_p0_93_port, Z(92) => state_main_in_p0_92_port, 
               Z(91) => state_main_in_p0_91_port, Z(90) => 
               state_main_in_p0_90_port, Z(89) => state_main_in_p0_89_port, 
               Z(88) => state_main_in_p0_88_port, Z(87) => 
               state_main_in_p0_87_port, Z(86) => state_main_in_p0_86_port, 
               Z(85) => state_main_in_p0_85_port, Z(84) => 
               state_main_in_p0_84_port, Z(83) => state_main_in_p0_83_port, 
               Z(82) => state_main_in_p0_82_port, Z(81) => 
               state_main_in_p0_81_port, Z(80) => state_main_in_p0_80_port, 
               Z(79) => state_main_in_p0_79_port, Z(78) => 
               state_main_in_p0_78_port, Z(77) => state_main_in_p0_77_port, 
               Z(76) => state_main_in_p0_76_port, Z(75) => 
               state_main_in_p0_75_port, Z(74) => state_main_in_p0_74_port, 
               Z(73) => state_main_in_p0_73_port, Z(72) => 
               state_main_in_p0_72_port, Z(71) => state_main_in_p0_71_port, 
               Z(70) => state_main_in_p0_70_port, Z(69) => 
               state_main_in_p0_69_port, Z(68) => state_main_in_p0_68_port, 
               Z(67) => state_main_in_p0_67_port, Z(66) => 
               state_main_in_p0_66_port, Z(65) => state_main_in_p0_65_port, 
               Z(64) => state_main_in_p0_64_port, Z(63) => 
               state_main_in_p0_63_port, Z(62) => state_main_in_p0_62_port, 
               Z(61) => state_main_in_p0_61_port, Z(60) => 
               state_main_in_p0_60_port, Z(59) => state_main_in_p0_59_port, 
               Z(58) => state_main_in_p0_58_port, Z(57) => 
               state_main_in_p0_57_port, Z(56) => state_main_in_p0_56_port, 
               Z(55) => state_main_in_p0_55_port, Z(54) => 
               state_main_in_p0_54_port, Z(53) => state_main_in_p0_53_port, 
               Z(52) => state_main_in_p0_52_port, Z(51) => 
               state_main_in_p0_51_port, Z(50) => state_main_in_p0_50_port, 
               Z(49) => state_main_in_p0_49_port, Z(48) => 
               state_main_in_p0_48_port, Z(47) => state_main_in_p0_47_port, 
               Z(46) => state_main_in_p0_46_port, Z(45) => 
               state_main_in_p0_45_port, Z(44) => state_main_in_p0_44_port, 
               Z(43) => state_main_in_p0_43_port, Z(42) => 
               state_main_in_p0_42_port, Z(41) => state_main_in_p0_41_port, 
               Z(40) => state_main_in_p0_40_port, Z(39) => 
               state_main_in_p0_39_port, Z(38) => state_main_in_p0_38_port, 
               Z(37) => state_main_in_p0_37_port, Z(36) => 
               state_main_in_p0_36_port, Z(35) => state_main_in_p0_35_port, 
               Z(34) => state_main_in_p0_34_port, Z(33) => 
               state_main_in_p0_33_port, Z(32) => state_main_in_p0_32_port, 
               Z(31) => state_main_in_p0_31_port, Z(30) => 
               state_main_in_p0_30_port, Z(29) => state_main_in_p0_29_port, 
               Z(28) => state_main_in_p0_28_port, Z(27) => 
               state_main_in_p0_27_port, Z(26) => state_main_in_p0_26_port, 
               Z(25) => state_main_in_p0_25_port, Z(24) => 
               state_main_in_p0_24_port, Z(23) => state_main_in_p0_23_port, 
               Z(22) => state_main_in_p0_22_port, Z(21) => 
               state_main_in_p0_21_port, Z(20) => state_main_in_p0_20_port, 
               Z(19) => state_main_in_p0_19_port, Z(18) => 
               state_main_in_p0_18_port, Z(17) => state_main_in_p0_17_port, 
               Z(16) => state_main_in_p0_16_port, Z(15) => 
               state_main_in_p0_15_port, Z(14) => state_main_in_p0_14_port, 
               Z(13) => state_main_in_p0_13_port, Z(12) => 
               state_main_in_p0_12_port, Z(11) => state_main_in_p0_11_port, 
               Z(10) => state_main_in_p0_10_port, Z(9) => 
               state_main_in_p0_9_port, Z(8) => state_main_in_p0_8_port, Z(7) 
               => state_main_in_p0_7_port, Z(6) => state_main_in_p0_6_port, 
               Z(5) => state_main_in_p0_5_port, Z(4) => state_main_in_p0_4_port
               , Z(3) => state_main_in_p0_3_port, Z(2) => 
               state_main_in_p0_2_port, Z(1) => state_main_in_p0_1_port, Z(0) 
               => state_main_in_p0_0_port );
   B_22 : GTECH_BUF port map( A => N181, Z => N22);
   B_23 : GTECH_BUF port map( A => state_main_sel(1), Z => N23);
   C1646_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 128 )
      port map(
         -- Connections to port 'DATA1'
         DATA(127) => cyc_state_update_127_port, DATA(126) => 
               cyc_state_update_126_port, DATA(125) => 
               cyc_state_update_125_port, DATA(124) => 
               cyc_state_update_124_port, DATA(123) => 
               cyc_state_update_123_port, DATA(122) => 
               cyc_state_update_122_port, DATA(121) => 
               cyc_state_update_121_port, DATA(120) => 
               cyc_state_update_120_port, DATA(119) => 
               cyc_state_update_119_port, DATA(118) => 
               cyc_state_update_118_port, DATA(117) => 
               cyc_state_update_117_port, DATA(116) => 
               cyc_state_update_116_port, DATA(115) => 
               cyc_state_update_115_port, DATA(114) => 
               cyc_state_update_114_port, DATA(113) => 
               cyc_state_update_113_port, DATA(112) => 
               cyc_state_update_112_port, DATA(111) => 
               cyc_state_update_111_port, DATA(110) => 
               cyc_state_update_110_port, DATA(109) => 
               cyc_state_update_109_port, DATA(108) => 
               cyc_state_update_108_port, DATA(107) => 
               cyc_state_update_107_port, DATA(106) => 
               cyc_state_update_106_port, DATA(105) => 
               cyc_state_update_105_port, DATA(104) => 
               cyc_state_update_104_port, DATA(103) => 
               cyc_state_update_103_port, DATA(102) => 
               cyc_state_update_102_port, DATA(101) => 
               cyc_state_update_101_port, DATA(100) => 
               cyc_state_update_100_port, DATA(99) => cyc_state_update_99_port,
               DATA(98) => cyc_state_update_98_port, DATA(97) => 
               cyc_state_update_97_port, DATA(96) => cyc_state_update_96_port, 
               DATA(95) => cyc_state_update_95_port, DATA(94) => 
               cyc_state_update_94_port, DATA(93) => cyc_state_update_93_port, 
               DATA(92) => cyc_state_update_92_port, DATA(91) => 
               cyc_state_update_91_port, DATA(90) => cyc_state_update_90_port, 
               DATA(89) => cyc_state_update_89_port, DATA(88) => 
               cyc_state_update_88_port, DATA(87) => cyc_state_update_87_port, 
               DATA(86) => cyc_state_update_86_port, DATA(85) => 
               cyc_state_update_85_port, DATA(84) => cyc_state_update_84_port, 
               DATA(83) => cyc_state_update_83_port, DATA(82) => 
               cyc_state_update_82_port, DATA(81) => cyc_state_update_81_port, 
               DATA(80) => cyc_state_update_80_port, DATA(79) => 
               cyc_state_update_79_port, DATA(78) => cyc_state_update_78_port, 
               DATA(77) => cyc_state_update_77_port, DATA(76) => 
               cyc_state_update_76_port, DATA(75) => cyc_state_update_75_port, 
               DATA(74) => cyc_state_update_74_port, DATA(73) => 
               cyc_state_update_73_port, DATA(72) => cyc_state_update_72_port, 
               DATA(71) => cyc_state_update_71_port, DATA(70) => 
               cyc_state_update_70_port, DATA(69) => cyc_state_update_69_port, 
               DATA(68) => cyc_state_update_68_port, DATA(67) => 
               cyc_state_update_67_port, DATA(66) => cyc_state_update_66_port, 
               DATA(65) => cyc_state_update_65_port, DATA(64) => 
               cyc_state_update_64_port, DATA(63) => cyc_state_update_63_port, 
               DATA(62) => cyc_state_update_62_port, DATA(61) => 
               cyc_state_update_61_port, DATA(60) => cyc_state_update_60_port, 
               DATA(59) => cyc_state_update_59_port, DATA(58) => 
               cyc_state_update_58_port, DATA(57) => cyc_state_update_57_port, 
               DATA(56) => cyc_state_update_56_port, DATA(55) => 
               cyc_state_update_55_port, DATA(54) => cyc_state_update_54_port, 
               DATA(53) => cyc_state_update_53_port, DATA(52) => 
               cyc_state_update_52_port, DATA(51) => cyc_state_update_51_port, 
               DATA(50) => cyc_state_update_50_port, DATA(49) => 
               cyc_state_update_49_port, DATA(48) => cyc_state_update_48_port, 
               DATA(47) => cyc_state_update_47_port, DATA(46) => 
               cyc_state_update_46_port, DATA(45) => cyc_state_update_45_port, 
               DATA(44) => cyc_state_update_44_port, DATA(43) => 
               cyc_state_update_43_port, DATA(42) => cyc_state_update_42_port, 
               DATA(41) => cyc_state_update_41_port, DATA(40) => 
               cyc_state_update_40_port, DATA(39) => cyc_state_update_39_port, 
               DATA(38) => cyc_state_update_38_port, DATA(37) => 
               cyc_state_update_37_port, DATA(36) => cyc_state_update_36_port, 
               DATA(35) => cyc_state_update_35_port, DATA(34) => 
               cyc_state_update_34_port, DATA(33) => cyc_state_update_33_port, 
               DATA(32) => cyc_state_update_32_port, DATA(31) => 
               cyc_state_update_31_port, DATA(30) => cyc_state_update_30_port, 
               DATA(29) => cyc_state_update_29_port, DATA(28) => 
               cyc_state_update_28_port, DATA(27) => cyc_state_update_27_port, 
               DATA(26) => cyc_state_update_26_port, DATA(25) => 
               cyc_state_update_25_port, DATA(24) => cyc_state_update_24_port, 
               DATA(23) => cyc_state_update_23_port, DATA(22) => 
               cyc_state_update_22_port, DATA(21) => cyc_state_update_21_port, 
               DATA(20) => cyc_state_update_20_port, DATA(19) => 
               cyc_state_update_19_port, DATA(18) => cyc_state_update_18_port, 
               DATA(17) => cyc_state_update_17_port, DATA(16) => 
               cyc_state_update_16_port, DATA(15) => cyc_state_update_15_port, 
               DATA(14) => cyc_state_update_14_port, DATA(13) => 
               cyc_state_update_13_port, DATA(12) => cyc_state_update_12_port, 
               DATA(11) => cyc_state_update_11_port, DATA(10) => 
               cyc_state_update_10_port, DATA(9) => cyc_state_update_9_port, 
               DATA(8) => cyc_state_update_8_port, DATA(7) => 
               cyc_state_update_7_port, DATA(6) => cyc_state_update_6_port, 
               DATA(5) => cyc_state_update_5_port, DATA(4) => 
               cyc_state_update_4_port, DATA(3) => cyc_state_update_3_port, 
               DATA(2) => cyc_state_update_2_port, DATA(1) => 
               cyc_state_update_1_port, DATA(0) => cyc_state_update_0_port, 
         -- Connections to port 'DATA2'
         DATA(255) => perm_output_255_port, DATA(254) => perm_output_254_port, 
               DATA(253) => perm_output_253_port, DATA(252) => 
               perm_output_252_port, DATA(251) => perm_output_251_port, 
               DATA(250) => perm_output_250_port, DATA(249) => 
               perm_output_249_port, DATA(248) => perm_output_248_port, 
               DATA(247) => perm_output_247_port, DATA(246) => 
               perm_output_246_port, DATA(245) => perm_output_245_port, 
               DATA(244) => perm_output_244_port, DATA(243) => 
               perm_output_243_port, DATA(242) => perm_output_242_port, 
               DATA(241) => perm_output_241_port, DATA(240) => 
               perm_output_240_port, DATA(239) => perm_output_239_port, 
               DATA(238) => perm_output_238_port, DATA(237) => 
               perm_output_237_port, DATA(236) => perm_output_236_port, 
               DATA(235) => perm_output_235_port, DATA(234) => 
               perm_output_234_port, DATA(233) => perm_output_233_port, 
               DATA(232) => perm_output_232_port, DATA(231) => 
               perm_output_231_port, DATA(230) => perm_output_230_port, 
               DATA(229) => perm_output_229_port, DATA(228) => 
               perm_output_228_port, DATA(227) => perm_output_227_port, 
               DATA(226) => perm_output_226_port, DATA(225) => 
               perm_output_225_port, DATA(224) => perm_output_224_port, 
               DATA(223) => perm_output_223_port, DATA(222) => 
               perm_output_222_port, DATA(221) => perm_output_221_port, 
               DATA(220) => perm_output_220_port, DATA(219) => 
               perm_output_219_port, DATA(218) => perm_output_218_port, 
               DATA(217) => perm_output_217_port, DATA(216) => 
               perm_output_216_port, DATA(215) => perm_output_215_port, 
               DATA(214) => perm_output_214_port, DATA(213) => 
               perm_output_213_port, DATA(212) => perm_output_212_port, 
               DATA(211) => perm_output_211_port, DATA(210) => 
               perm_output_210_port, DATA(209) => perm_output_209_port, 
               DATA(208) => perm_output_208_port, DATA(207) => 
               perm_output_207_port, DATA(206) => perm_output_206_port, 
               DATA(205) => perm_output_205_port, DATA(204) => 
               perm_output_204_port, DATA(203) => perm_output_203_port, 
               DATA(202) => perm_output_202_port, DATA(201) => 
               perm_output_201_port, DATA(200) => perm_output_200_port, 
               DATA(199) => perm_output_199_port, DATA(198) => 
               perm_output_198_port, DATA(197) => perm_output_197_port, 
               DATA(196) => perm_output_196_port, DATA(195) => 
               perm_output_195_port, DATA(194) => perm_output_194_port, 
               DATA(193) => perm_output_193_port, DATA(192) => 
               perm_output_192_port, DATA(191) => perm_output_191_port, 
               DATA(190) => perm_output_190_port, DATA(189) => 
               perm_output_189_port, DATA(188) => perm_output_188_port, 
               DATA(187) => perm_output_187_port, DATA(186) => 
               perm_output_186_port, DATA(185) => perm_output_185_port, 
               DATA(184) => perm_output_184_port, DATA(183) => 
               perm_output_183_port, DATA(182) => perm_output_182_port, 
               DATA(181) => perm_output_181_port, DATA(180) => 
               perm_output_180_port, DATA(179) => perm_output_179_port, 
               DATA(178) => perm_output_178_port, DATA(177) => 
               perm_output_177_port, DATA(176) => perm_output_176_port, 
               DATA(175) => perm_output_175_port, DATA(174) => 
               perm_output_174_port, DATA(173) => perm_output_173_port, 
               DATA(172) => perm_output_172_port, DATA(171) => 
               perm_output_171_port, DATA(170) => perm_output_170_port, 
               DATA(169) => perm_output_169_port, DATA(168) => 
               perm_output_168_port, DATA(167) => perm_output_167_port, 
               DATA(166) => perm_output_166_port, DATA(165) => 
               perm_output_165_port, DATA(164) => perm_output_164_port, 
               DATA(163) => perm_output_163_port, DATA(162) => 
               perm_output_162_port, DATA(161) => perm_output_161_port, 
               DATA(160) => perm_output_160_port, DATA(159) => 
               perm_output_159_port, DATA(158) => perm_output_158_port, 
               DATA(157) => perm_output_157_port, DATA(156) => 
               perm_output_156_port, DATA(155) => perm_output_155_port, 
               DATA(154) => perm_output_154_port, DATA(153) => 
               perm_output_153_port, DATA(152) => perm_output_152_port, 
               DATA(151) => perm_output_151_port, DATA(150) => 
               perm_output_150_port, DATA(149) => perm_output_149_port, 
               DATA(148) => perm_output_148_port, DATA(147) => 
               perm_output_147_port, DATA(146) => perm_output_146_port, 
               DATA(145) => perm_output_145_port, DATA(144) => 
               perm_output_144_port, DATA(143) => perm_output_143_port, 
               DATA(142) => perm_output_142_port, DATA(141) => 
               perm_output_141_port, DATA(140) => perm_output_140_port, 
               DATA(139) => perm_output_139_port, DATA(138) => 
               perm_output_138_port, DATA(137) => perm_output_137_port, 
               DATA(136) => perm_output_136_port, DATA(135) => 
               perm_output_135_port, DATA(134) => perm_output_134_port, 
               DATA(133) => perm_output_133_port, DATA(132) => 
               perm_output_132_port, DATA(131) => perm_output_131_port, 
               DATA(130) => perm_output_130_port, DATA(129) => 
               perm_output_129_port, DATA(128) => perm_output_128_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N24, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N25, 
         -- Connections to port 'Z'
         Z(127) => N440, Z(126) => N439, Z(125) => N438, Z(124) => N437, Z(123)
               => N436, Z(122) => N435, Z(121) => N434, Z(120) => N433, Z(119) 
               => N432, Z(118) => N431, Z(117) => N430, Z(116) => N429, Z(115) 
               => N428, Z(114) => N427, Z(113) => N426, Z(112) => N425, Z(111) 
               => N424, Z(110) => N423, Z(109) => N422, Z(108) => N421, Z(107) 
               => N420, Z(106) => N419, Z(105) => N418, Z(104) => N417, Z(103) 
               => N416, Z(102) => N415, Z(101) => N414, Z(100) => N413, Z(99) 
               => N412, Z(98) => N411, Z(97) => N410, Z(96) => N409, Z(95) => 
               N408, Z(94) => N407, Z(93) => N406, Z(92) => N405, Z(91) => N404
               , Z(90) => N403, Z(89) => N402, Z(88) => N401, Z(87) => N400, 
               Z(86) => N399, Z(85) => N398, Z(84) => N397, Z(83) => N396, 
               Z(82) => N395, Z(81) => N394, Z(80) => N393, Z(79) => N392, 
               Z(78) => N391, Z(77) => N390, Z(76) => N389, Z(75) => N388, 
               Z(74) => N387, Z(73) => N386, Z(72) => N385, Z(71) => N384, 
               Z(70) => N383, Z(69) => N382, Z(68) => N381, Z(67) => N380, 
               Z(66) => N379, Z(65) => N378, Z(64) => N377, Z(63) => N376, 
               Z(62) => N375, Z(61) => N374, Z(60) => N373, Z(59) => N372, 
               Z(58) => N371, Z(57) => N370, Z(56) => N369, Z(55) => N368, 
               Z(54) => N367, Z(53) => N366, Z(52) => N365, Z(51) => N364, 
               Z(50) => N363, Z(49) => N362, Z(48) => N361, Z(47) => N360, 
               Z(46) => N359, Z(45) => N358, Z(44) => N357, Z(43) => N356, 
               Z(42) => N355, Z(41) => N354, Z(40) => N353, Z(39) => N352, 
               Z(38) => N351, Z(37) => N350, Z(36) => N349, Z(35) => N348, 
               Z(34) => N347, Z(33) => N346, Z(32) => N345, Z(31) => N344, 
               Z(30) => N343, Z(29) => N342, Z(28) => N341, Z(27) => N340, 
               Z(26) => N339, Z(25) => N338, Z(24) => N337, Z(23) => N336, 
               Z(22) => N335, Z(21) => N334, Z(20) => N333, Z(19) => N332, 
               Z(18) => N331, Z(17) => N330, Z(16) => N329, Z(15) => N328, 
               Z(14) => N327, Z(13) => N326, Z(12) => N325, Z(11) => N324, 
               Z(10) => N323, Z(9) => N322, Z(8) => N321, Z(7) => N320, Z(6) =>
               N319, Z(5) => N318, Z(4) => N317, Z(3) => N316, Z(2) => N315, 
               Z(1) => N314, Z(0) => N313 );
   B_24 : GTECH_BUF port map( A => N312, Z => N24);
   B_25 : GTECH_BUF port map( A => state_main_sel(2), Z => N25);
   C1647_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 128 )
      port map(
         -- Connections to port 'DATA1'
         DATA(127) => N440, DATA(126) => N439, DATA(125) => N438, DATA(124) => 
               N437, DATA(123) => N436, DATA(122) => N435, DATA(121) => N434, 
               DATA(120) => N433, DATA(119) => N432, DATA(118) => N431, 
               DATA(117) => N430, DATA(116) => N429, DATA(115) => N428, 
               DATA(114) => N427, DATA(113) => N426, DATA(112) => N425, 
               DATA(111) => N424, DATA(110) => N423, DATA(109) => N422, 
               DATA(108) => N421, DATA(107) => N420, DATA(106) => N419, 
               DATA(105) => N418, DATA(104) => N417, DATA(103) => N416, 
               DATA(102) => N415, DATA(101) => N414, DATA(100) => N413, 
               DATA(99) => N412, DATA(98) => N411, DATA(97) => N410, DATA(96) 
               => N409, DATA(95) => N408, DATA(94) => N407, DATA(93) => N406, 
               DATA(92) => N405, DATA(91) => N404, DATA(90) => N403, DATA(89) 
               => N402, DATA(88) => N401, DATA(87) => N400, DATA(86) => N399, 
               DATA(85) => N398, DATA(84) => N397, DATA(83) => N396, DATA(82) 
               => N395, DATA(81) => N394, DATA(80) => N393, DATA(79) => N392, 
               DATA(78) => N391, DATA(77) => N390, DATA(76) => N389, DATA(75) 
               => N388, DATA(74) => N387, DATA(73) => N386, DATA(72) => N385, 
               DATA(71) => N384, DATA(70) => N383, DATA(69) => N382, DATA(68) 
               => N381, DATA(67) => N380, DATA(66) => N379, DATA(65) => N378, 
               DATA(64) => N377, DATA(63) => N376, DATA(62) => N375, DATA(61) 
               => N374, DATA(60) => N373, DATA(59) => N372, DATA(58) => N371, 
               DATA(57) => N370, DATA(56) => N369, DATA(55) => N368, DATA(54) 
               => N367, DATA(53) => N366, DATA(52) => N365, DATA(51) => N364, 
               DATA(50) => N363, DATA(49) => N362, DATA(48) => N361, DATA(47) 
               => N360, DATA(46) => N359, DATA(45) => N358, DATA(44) => N357, 
               DATA(43) => N356, DATA(42) => N355, DATA(41) => N354, DATA(40) 
               => N353, DATA(39) => N352, DATA(38) => N351, DATA(37) => N350, 
               DATA(36) => N349, DATA(35) => N348, DATA(34) => N347, DATA(33) 
               => N346, DATA(32) => N345, DATA(31) => N344, DATA(30) => N343, 
               DATA(29) => N342, DATA(28) => N341, DATA(27) => N340, DATA(26) 
               => N339, DATA(25) => N338, DATA(24) => N337, DATA(23) => N336, 
               DATA(22) => N335, DATA(21) => N334, DATA(20) => N333, DATA(19) 
               => N332, DATA(18) => N331, DATA(17) => N330, DATA(16) => N329, 
               DATA(15) => N328, DATA(14) => N327, DATA(13) => N326, DATA(12) 
               => N325, DATA(11) => N324, DATA(10) => N323, DATA(9) => N322, 
               DATA(8) => N321, DATA(7) => N320, DATA(6) => N319, DATA(5) => 
               N318, DATA(4) => N317, DATA(3) => N316, DATA(2) => N315, DATA(1)
               => N314, DATA(0) => N313, 
         -- Connections to port 'DATA2'
         DATA(255) => X_Logic0_port, DATA(254) => X_Logic0_port, DATA(253) => 
               X_Logic0_port, DATA(252) => X_Logic0_port, DATA(251) => 
               X_Logic0_port, DATA(250) => X_Logic0_port, DATA(249) => 
               X_Logic0_port, DATA(248) => X_Logic0_port, DATA(247) => 
               X_Logic0_port, DATA(246) => X_Logic0_port, DATA(245) => 
               X_Logic0_port, DATA(244) => X_Logic0_port, DATA(243) => 
               X_Logic0_port, DATA(242) => X_Logic0_port, DATA(241) => 
               X_Logic0_port, DATA(240) => X_Logic0_port, DATA(239) => 
               X_Logic0_port, DATA(238) => X_Logic0_port, DATA(237) => 
               X_Logic0_port, DATA(236) => X_Logic0_port, DATA(235) => 
               X_Logic0_port, DATA(234) => X_Logic0_port, DATA(233) => 
               X_Logic0_port, DATA(232) => X_Logic0_port, DATA(231) => 
               X_Logic0_port, DATA(230) => X_Logic0_port, DATA(229) => 
               X_Logic0_port, DATA(228) => X_Logic0_port, DATA(227) => 
               X_Logic0_port, DATA(226) => X_Logic0_port, DATA(225) => 
               X_Logic0_port, DATA(224) => X_Logic0_port, DATA(223) => 
               X_Logic0_port, DATA(222) => X_Logic0_port, DATA(221) => 
               X_Logic0_port, DATA(220) => X_Logic0_port, DATA(219) => 
               X_Logic0_port, DATA(218) => X_Logic0_port, DATA(217) => 
               X_Logic0_port, DATA(216) => X_Logic0_port, DATA(215) => 
               X_Logic0_port, DATA(214) => X_Logic0_port, DATA(213) => 
               X_Logic0_port, DATA(212) => X_Logic0_port, DATA(211) => 
               X_Logic0_port, DATA(210) => X_Logic0_port, DATA(209) => 
               X_Logic0_port, DATA(208) => X_Logic0_port, DATA(207) => 
               X_Logic0_port, DATA(206) => X_Logic0_port, DATA(205) => 
               X_Logic0_port, DATA(204) => X_Logic0_port, DATA(203) => 
               X_Logic0_port, DATA(202) => X_Logic0_port, DATA(201) => 
               X_Logic0_port, DATA(200) => X_Logic0_port, DATA(199) => 
               X_Logic0_port, DATA(198) => X_Logic0_port, DATA(197) => 
               X_Logic0_port, DATA(196) => X_Logic0_port, DATA(195) => 
               X_Logic0_port, DATA(194) => X_Logic0_port, DATA(193) => 
               X_Logic0_port, DATA(192) => X_Logic0_port, DATA(191) => 
               X_Logic0_port, DATA(190) => X_Logic0_port, DATA(189) => 
               X_Logic0_port, DATA(188) => X_Logic0_port, DATA(187) => 
               X_Logic0_port, DATA(186) => X_Logic0_port, DATA(185) => 
               X_Logic0_port, DATA(184) => X_Logic0_port, DATA(183) => 
               X_Logic0_port, DATA(182) => X_Logic0_port, DATA(181) => 
               X_Logic0_port, DATA(180) => X_Logic0_port, DATA(179) => 
               X_Logic0_port, DATA(178) => X_Logic0_port, DATA(177) => 
               X_Logic0_port, DATA(176) => X_Logic0_port, DATA(175) => 
               X_Logic0_port, DATA(174) => X_Logic0_port, DATA(173) => 
               X_Logic0_port, DATA(172) => X_Logic0_port, DATA(171) => 
               X_Logic0_port, DATA(170) => X_Logic0_port, DATA(169) => 
               X_Logic0_port, DATA(168) => X_Logic0_port, DATA(167) => 
               X_Logic0_port, DATA(166) => X_Logic0_port, DATA(165) => 
               X_Logic0_port, DATA(164) => X_Logic0_port, DATA(163) => 
               X_Logic0_port, DATA(162) => X_Logic0_port, DATA(161) => 
               X_Logic0_port, DATA(160) => X_Logic0_port, DATA(159) => 
               X_Logic0_port, DATA(158) => X_Logic0_port, DATA(157) => 
               X_Logic0_port, DATA(156) => X_Logic0_port, DATA(155) => 
               X_Logic0_port, DATA(154) => X_Logic0_port, DATA(153) => 
               X_Logic0_port, DATA(152) => X_Logic0_port, DATA(151) => 
               X_Logic0_port, DATA(150) => X_Logic0_port, DATA(149) => 
               X_Logic0_port, DATA(148) => X_Logic0_port, DATA(147) => 
               X_Logic0_port, DATA(146) => X_Logic0_port, DATA(145) => 
               X_Logic0_port, DATA(144) => X_Logic0_port, DATA(143) => 
               X_Logic0_port, DATA(142) => X_Logic0_port, DATA(141) => 
               X_Logic0_port, DATA(140) => X_Logic0_port, DATA(139) => 
               X_Logic0_port, DATA(138) => X_Logic0_port, DATA(137) => 
               X_Logic0_port, DATA(136) => X_Logic0_port, DATA(135) => 
               X_Logic0_port, DATA(134) => X_Logic0_port, DATA(133) => 
               X_Logic0_port, DATA(132) => X_Logic0_port, DATA(131) => 
               X_Logic0_port, DATA(130) => X_Logic0_port, DATA(129) => 
               X_Logic0_port, DATA(128) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N26, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N27, 
         -- Connections to port 'Z'
         Z(127) => state_main_in_p1_127_port, Z(126) => 
               state_main_in_p1_126_port, Z(125) => state_main_in_p1_125_port, 
               Z(124) => state_main_in_p1_124_port, Z(123) => 
               state_main_in_p1_123_port, Z(122) => state_main_in_p1_122_port, 
               Z(121) => state_main_in_p1_121_port, Z(120) => 
               state_main_in_p1_120_port, Z(119) => state_main_in_p1_119_port, 
               Z(118) => state_main_in_p1_118_port, Z(117) => 
               state_main_in_p1_117_port, Z(116) => state_main_in_p1_116_port, 
               Z(115) => state_main_in_p1_115_port, Z(114) => 
               state_main_in_p1_114_port, Z(113) => state_main_in_p1_113_port, 
               Z(112) => state_main_in_p1_112_port, Z(111) => 
               state_main_in_p1_111_port, Z(110) => state_main_in_p1_110_port, 
               Z(109) => state_main_in_p1_109_port, Z(108) => 
               state_main_in_p1_108_port, Z(107) => state_main_in_p1_107_port, 
               Z(106) => state_main_in_p1_106_port, Z(105) => 
               state_main_in_p1_105_port, Z(104) => state_main_in_p1_104_port, 
               Z(103) => state_main_in_p1_103_port, Z(102) => 
               state_main_in_p1_102_port, Z(101) => state_main_in_p1_101_port, 
               Z(100) => state_main_in_p1_100_port, Z(99) => 
               state_main_in_p1_99_port, Z(98) => state_main_in_p1_98_port, 
               Z(97) => state_main_in_p1_97_port, Z(96) => 
               state_main_in_p1_96_port, Z(95) => state_main_in_p1_95_port, 
               Z(94) => state_main_in_p1_94_port, Z(93) => 
               state_main_in_p1_93_port, Z(92) => state_main_in_p1_92_port, 
               Z(91) => state_main_in_p1_91_port, Z(90) => 
               state_main_in_p1_90_port, Z(89) => state_main_in_p1_89_port, 
               Z(88) => state_main_in_p1_88_port, Z(87) => 
               state_main_in_p1_87_port, Z(86) => state_main_in_p1_86_port, 
               Z(85) => state_main_in_p1_85_port, Z(84) => 
               state_main_in_p1_84_port, Z(83) => state_main_in_p1_83_port, 
               Z(82) => state_main_in_p1_82_port, Z(81) => 
               state_main_in_p1_81_port, Z(80) => state_main_in_p1_80_port, 
               Z(79) => state_main_in_p1_79_port, Z(78) => 
               state_main_in_p1_78_port, Z(77) => state_main_in_p1_77_port, 
               Z(76) => state_main_in_p1_76_port, Z(75) => 
               state_main_in_p1_75_port, Z(74) => state_main_in_p1_74_port, 
               Z(73) => state_main_in_p1_73_port, Z(72) => 
               state_main_in_p1_72_port, Z(71) => state_main_in_p1_71_port, 
               Z(70) => state_main_in_p1_70_port, Z(69) => 
               state_main_in_p1_69_port, Z(68) => state_main_in_p1_68_port, 
               Z(67) => state_main_in_p1_67_port, Z(66) => 
               state_main_in_p1_66_port, Z(65) => state_main_in_p1_65_port, 
               Z(64) => state_main_in_p1_64_port, Z(63) => 
               state_main_in_p1_63_port, Z(62) => state_main_in_p1_62_port, 
               Z(61) => state_main_in_p1_61_port, Z(60) => 
               state_main_in_p1_60_port, Z(59) => state_main_in_p1_59_port, 
               Z(58) => state_main_in_p1_58_port, Z(57) => 
               state_main_in_p1_57_port, Z(56) => state_main_in_p1_56_port, 
               Z(55) => state_main_in_p1_55_port, Z(54) => 
               state_main_in_p1_54_port, Z(53) => state_main_in_p1_53_port, 
               Z(52) => state_main_in_p1_52_port, Z(51) => 
               state_main_in_p1_51_port, Z(50) => state_main_in_p1_50_port, 
               Z(49) => state_main_in_p1_49_port, Z(48) => 
               state_main_in_p1_48_port, Z(47) => state_main_in_p1_47_port, 
               Z(46) => state_main_in_p1_46_port, Z(45) => 
               state_main_in_p1_45_port, Z(44) => state_main_in_p1_44_port, 
               Z(43) => state_main_in_p1_43_port, Z(42) => 
               state_main_in_p1_42_port, Z(41) => state_main_in_p1_41_port, 
               Z(40) => state_main_in_p1_40_port, Z(39) => 
               state_main_in_p1_39_port, Z(38) => state_main_in_p1_38_port, 
               Z(37) => state_main_in_p1_37_port, Z(36) => 
               state_main_in_p1_36_port, Z(35) => state_main_in_p1_35_port, 
               Z(34) => state_main_in_p1_34_port, Z(33) => 
               state_main_in_p1_33_port, Z(32) => state_main_in_p1_32_port, 
               Z(31) => state_main_in_p1_31_port, Z(30) => 
               state_main_in_p1_30_port, Z(29) => state_main_in_p1_29_port, 
               Z(28) => state_main_in_p1_28_port, Z(27) => 
               state_main_in_p1_27_port, Z(26) => state_main_in_p1_26_port, 
               Z(25) => state_main_in_p1_25_port, Z(24) => 
               state_main_in_p1_24_port, Z(23) => state_main_in_p1_23_port, 
               Z(22) => state_main_in_p1_22_port, Z(21) => 
               state_main_in_p1_21_port, Z(20) => state_main_in_p1_20_port, 
               Z(19) => state_main_in_p1_19_port, Z(18) => 
               state_main_in_p1_18_port, Z(17) => state_main_in_p1_17_port, 
               Z(16) => state_main_in_p1_16_port, Z(15) => 
               state_main_in_p1_15_port, Z(14) => state_main_in_p1_14_port, 
               Z(13) => state_main_in_p1_13_port, Z(12) => 
               state_main_in_p1_12_port, Z(11) => state_main_in_p1_11_port, 
               Z(10) => state_main_in_p1_10_port, Z(9) => 
               state_main_in_p1_9_port, Z(8) => state_main_in_p1_8_port, Z(7) 
               => state_main_in_p1_7_port, Z(6) => state_main_in_p1_6_port, 
               Z(5) => state_main_in_p1_5_port, Z(4) => state_main_in_p1_4_port
               , Z(3) => state_main_in_p1_3_port, Z(2) => 
               state_main_in_p1_2_port, Z(1) => state_main_in_p1_1_port, Z(0) 
               => state_main_in_p1_0_port );
   B_26 : GTECH_BUF port map( A => N311, Z => N26);
   B_27 : GTECH_BUF port map( A => state_main_sel(3), Z => N27);
   C1648_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 128 )
      port map(
         -- Connections to port 'DATA1'
         DATA(127) => plane_2_input_127_port, DATA(126) => 
               plane_2_input_126_port, DATA(125) => plane_2_input_125_port, 
               DATA(124) => plane_2_input_124_port, DATA(123) => 
               plane_2_input_123_port, DATA(122) => plane_2_input_122_port, 
               DATA(121) => plane_2_input_121_port, DATA(120) => 
               plane_2_input_120_port, DATA(119) => plane_2_input_119_port, 
               DATA(118) => plane_2_input_118_port, DATA(117) => 
               plane_2_input_117_port, DATA(116) => plane_2_input_116_port, 
               DATA(115) => plane_2_input_115_port, DATA(114) => 
               plane_2_input_114_port, DATA(113) => plane_2_input_113_port, 
               DATA(112) => plane_2_input_112_port, DATA(111) => 
               plane_2_input_111_port, DATA(110) => plane_2_input_110_port, 
               DATA(109) => plane_2_input_109_port, DATA(108) => 
               plane_2_input_108_port, DATA(107) => plane_2_input_107_port, 
               DATA(106) => plane_2_input_106_port, DATA(105) => 
               plane_2_input_105_port, DATA(104) => plane_2_input_104_port, 
               DATA(103) => plane_2_input_103_port, DATA(102) => 
               plane_2_input_102_port, DATA(101) => plane_2_input_101_port, 
               DATA(100) => plane_2_input_100_port, DATA(99) => 
               plane_2_input_99_port, DATA(98) => plane_2_input_98_port, 
               DATA(97) => plane_2_input_97_port, DATA(96) => 
               plane_2_input_96_port, DATA(95) => plane_2_input_95_port, 
               DATA(94) => plane_2_input_94_port, DATA(93) => 
               plane_2_input_93_port, DATA(92) => plane_2_input_92_port, 
               DATA(91) => plane_2_input_91_port, DATA(90) => 
               plane_2_input_90_port, DATA(89) => plane_2_input_89_port, 
               DATA(88) => plane_2_input_88_port, DATA(87) => 
               plane_2_input_87_port, DATA(86) => plane_2_input_86_port, 
               DATA(85) => plane_2_input_85_port, DATA(84) => 
               plane_2_input_84_port, DATA(83) => plane_2_input_83_port, 
               DATA(82) => plane_2_input_82_port, DATA(81) => 
               plane_2_input_81_port, DATA(80) => plane_2_input_80_port, 
               DATA(79) => plane_2_input_79_port, DATA(78) => 
               plane_2_input_78_port, DATA(77) => plane_2_input_77_port, 
               DATA(76) => plane_2_input_76_port, DATA(75) => 
               plane_2_input_75_port, DATA(74) => plane_2_input_74_port, 
               DATA(73) => plane_2_input_73_port, DATA(72) => 
               plane_2_input_72_port, DATA(71) => plane_2_input_71_port, 
               DATA(70) => plane_2_input_70_port, DATA(69) => 
               plane_2_input_69_port, DATA(68) => plane_2_input_68_port, 
               DATA(67) => plane_2_input_67_port, DATA(66) => 
               plane_2_input_66_port, DATA(65) => plane_2_input_65_port, 
               DATA(64) => plane_2_input_64_port, DATA(63) => 
               plane_2_input_63_port, DATA(62) => plane_2_input_62_port, 
               DATA(61) => plane_2_input_61_port, DATA(60) => 
               plane_2_input_60_port, DATA(59) => plane_2_input_59_port, 
               DATA(58) => plane_2_input_58_port, DATA(57) => 
               plane_2_input_57_port, DATA(56) => plane_2_input_56_port, 
               DATA(55) => plane_2_input_55_port, DATA(54) => 
               plane_2_input_54_port, DATA(53) => plane_2_input_53_port, 
               DATA(52) => plane_2_input_52_port, DATA(51) => 
               plane_2_input_51_port, DATA(50) => plane_2_input_50_port, 
               DATA(49) => plane_2_input_49_port, DATA(48) => 
               plane_2_input_48_port, DATA(47) => plane_2_input_47_port, 
               DATA(46) => plane_2_input_46_port, DATA(45) => 
               plane_2_input_45_port, DATA(44) => plane_2_input_44_port, 
               DATA(43) => plane_2_input_43_port, DATA(42) => 
               plane_2_input_42_port, DATA(41) => plane_2_input_41_port, 
               DATA(40) => plane_2_input_40_port, DATA(39) => 
               plane_2_input_39_port, DATA(38) => plane_2_input_38_port, 
               DATA(37) => plane_2_input_37_port, DATA(36) => 
               plane_2_input_36_port, DATA(35) => plane_2_input_35_port, 
               DATA(34) => plane_2_input_34_port, DATA(33) => 
               plane_2_input_33_port, DATA(32) => plane_2_input_32_port, 
               DATA(31) => fb_prime_7_port, DATA(30) => fb_prime_6_port, 
               DATA(29) => fb_prime_5_port, DATA(28) => fb_prime_4_port, 
               DATA(27) => fb_prime_3_port, DATA(26) => fb_prime_2_port, 
               DATA(25) => fb_prime_1_port, DATA(24) => fb_prime_0_port, 
               DATA(23) => plane_2_input_23, DATA(22) => plane_2_input_22, 
               DATA(21) => plane_2_input_21, DATA(20) => plane_2_input_20, 
               DATA(19) => plane_2_input_19, DATA(18) => plane_2_input_18, 
               DATA(17) => plane_2_input_17, DATA(16) => plane_2_input_16, 
               DATA(15) => plane_2_input_15, DATA(14) => plane_2_input_14, 
               DATA(13) => plane_2_input_13, DATA(12) => plane_2_input_12, 
               DATA(11) => plane_2_input_11, DATA(10) => plane_2_input_10, 
               DATA(9) => plane_2_input_9, DATA(8) => plane_2_input_8, DATA(7) 
               => plane_2_input_7, DATA(6) => plane_2_input_6, DATA(5) => 
               plane_2_input_5, DATA(4) => plane_2_input_4, DATA(3) => 
               plane_2_input_3, DATA(2) => plane_2_input_2, DATA(1) => 
               plane_2_input_1, DATA(0) => plane_2_input_0, 
         -- Connections to port 'DATA2'
         DATA(255) => perm_output_383_port, DATA(254) => perm_output_382_port, 
               DATA(253) => perm_output_381_port, DATA(252) => 
               perm_output_380_port, DATA(251) => perm_output_379_port, 
               DATA(250) => perm_output_378_port, DATA(249) => 
               perm_output_377_port, DATA(248) => perm_output_376_port, 
               DATA(247) => perm_output_375_port, DATA(246) => 
               perm_output_374_port, DATA(245) => perm_output_373_port, 
               DATA(244) => perm_output_372_port, DATA(243) => 
               perm_output_371_port, DATA(242) => perm_output_370_port, 
               DATA(241) => perm_output_369_port, DATA(240) => 
               perm_output_368_port, DATA(239) => perm_output_367_port, 
               DATA(238) => perm_output_366_port, DATA(237) => 
               perm_output_365_port, DATA(236) => perm_output_364_port, 
               DATA(235) => perm_output_363_port, DATA(234) => 
               perm_output_362_port, DATA(233) => perm_output_361_port, 
               DATA(232) => perm_output_360_port, DATA(231) => 
               perm_output_359_port, DATA(230) => perm_output_358_port, 
               DATA(229) => perm_output_357_port, DATA(228) => 
               perm_output_356_port, DATA(227) => perm_output_355_port, 
               DATA(226) => perm_output_354_port, DATA(225) => 
               perm_output_353_port, DATA(224) => perm_output_352_port, 
               DATA(223) => perm_output_351_port, DATA(222) => 
               perm_output_350_port, DATA(221) => perm_output_349_port, 
               DATA(220) => perm_output_348_port, DATA(219) => 
               perm_output_347_port, DATA(218) => perm_output_346_port, 
               DATA(217) => perm_output_345_port, DATA(216) => 
               perm_output_344_port, DATA(215) => perm_output_343_port, 
               DATA(214) => perm_output_342_port, DATA(213) => 
               perm_output_341_port, DATA(212) => perm_output_340_port, 
               DATA(211) => perm_output_339_port, DATA(210) => 
               perm_output_338_port, DATA(209) => perm_output_337_port, 
               DATA(208) => perm_output_336_port, DATA(207) => 
               perm_output_335_port, DATA(206) => perm_output_334_port, 
               DATA(205) => perm_output_333_port, DATA(204) => 
               perm_output_332_port, DATA(203) => perm_output_331_port, 
               DATA(202) => perm_output_330_port, DATA(201) => 
               perm_output_329_port, DATA(200) => perm_output_328_port, 
               DATA(199) => perm_output_327_port, DATA(198) => 
               perm_output_326_port, DATA(197) => perm_output_325_port, 
               DATA(196) => perm_output_324_port, DATA(195) => 
               perm_output_323_port, DATA(194) => perm_output_322_port, 
               DATA(193) => perm_output_321_port, DATA(192) => 
               perm_output_320_port, DATA(191) => perm_output_319_port, 
               DATA(190) => perm_output_318_port, DATA(189) => 
               perm_output_317_port, DATA(188) => perm_output_316_port, 
               DATA(187) => perm_output_315_port, DATA(186) => 
               perm_output_314_port, DATA(185) => perm_output_313_port, 
               DATA(184) => perm_output_312_port, DATA(183) => 
               perm_output_311_port, DATA(182) => perm_output_310_port, 
               DATA(181) => perm_output_309_port, DATA(180) => 
               perm_output_308_port, DATA(179) => perm_output_307_port, 
               DATA(178) => perm_output_306_port, DATA(177) => 
               perm_output_305_port, DATA(176) => perm_output_304_port, 
               DATA(175) => perm_output_303_port, DATA(174) => 
               perm_output_302_port, DATA(173) => perm_output_301_port, 
               DATA(172) => perm_output_300_port, DATA(171) => 
               perm_output_299_port, DATA(170) => perm_output_298_port, 
               DATA(169) => perm_output_297_port, DATA(168) => 
               perm_output_296_port, DATA(167) => perm_output_295_port, 
               DATA(166) => perm_output_294_port, DATA(165) => 
               perm_output_293_port, DATA(164) => perm_output_292_port, 
               DATA(163) => perm_output_291_port, DATA(162) => 
               perm_output_290_port, DATA(161) => perm_output_289_port, 
               DATA(160) => perm_output_288_port, DATA(159) => 
               perm_output_287_port, DATA(158) => perm_output_286_port, 
               DATA(157) => perm_output_285_port, DATA(156) => 
               perm_output_284_port, DATA(155) => perm_output_283_port, 
               DATA(154) => perm_output_282_port, DATA(153) => 
               perm_output_281_port, DATA(152) => perm_output_280_port, 
               DATA(151) => perm_output_279_port, DATA(150) => 
               perm_output_278_port, DATA(149) => perm_output_277_port, 
               DATA(148) => perm_output_276_port, DATA(147) => 
               perm_output_275_port, DATA(146) => perm_output_274_port, 
               DATA(145) => perm_output_273_port, DATA(144) => 
               perm_output_272_port, DATA(143) => perm_output_271_port, 
               DATA(142) => perm_output_270_port, DATA(141) => 
               perm_output_269_port, DATA(140) => perm_output_268_port, 
               DATA(139) => perm_output_267_port, DATA(138) => 
               perm_output_266_port, DATA(137) => perm_output_265_port, 
               DATA(136) => perm_output_264_port, DATA(135) => 
               perm_output_263_port, DATA(134) => perm_output_262_port, 
               DATA(133) => perm_output_261_port, DATA(132) => 
               perm_output_260_port, DATA(131) => perm_output_259_port, 
               DATA(130) => perm_output_258_port, DATA(129) => 
               perm_output_257_port, DATA(128) => perm_output_256_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N28, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N29, 
         -- Connections to port 'Z'
         Z(127) => N570, Z(126) => N569, Z(125) => N568, Z(124) => N567, Z(123)
               => N566, Z(122) => N565, Z(121) => N564, Z(120) => N563, Z(119) 
               => N562, Z(118) => N561, Z(117) => N560, Z(116) => N559, Z(115) 
               => N558, Z(114) => N557, Z(113) => N556, Z(112) => N555, Z(111) 
               => N554, Z(110) => N553, Z(109) => N552, Z(108) => N551, Z(107) 
               => N550, Z(106) => N549, Z(105) => N548, Z(104) => N547, Z(103) 
               => N546, Z(102) => N545, Z(101) => N544, Z(100) => N543, Z(99) 
               => N542, Z(98) => N541, Z(97) => N540, Z(96) => N539, Z(95) => 
               N538, Z(94) => N537, Z(93) => N536, Z(92) => N535, Z(91) => N534
               , Z(90) => N533, Z(89) => N532, Z(88) => N531, Z(87) => N530, 
               Z(86) => N529, Z(85) => N528, Z(84) => N527, Z(83) => N526, 
               Z(82) => N525, Z(81) => N524, Z(80) => N523, Z(79) => N522, 
               Z(78) => N521, Z(77) => N520, Z(76) => N519, Z(75) => N518, 
               Z(74) => N517, Z(73) => N516, Z(72) => N515, Z(71) => N514, 
               Z(70) => N513, Z(69) => N512, Z(68) => N511, Z(67) => N510, 
               Z(66) => N509, Z(65) => N508, Z(64) => N507, Z(63) => N506, 
               Z(62) => N505, Z(61) => N504, Z(60) => N503, Z(59) => N502, 
               Z(58) => N501, Z(57) => N500, Z(56) => N499, Z(55) => N498, 
               Z(54) => N497, Z(53) => N496, Z(52) => N495, Z(51) => N494, 
               Z(50) => N493, Z(49) => N492, Z(48) => N491, Z(47) => N490, 
               Z(46) => N489, Z(45) => N488, Z(44) => N487, Z(43) => N486, 
               Z(42) => N485, Z(41) => N484, Z(40) => N483, Z(39) => N482, 
               Z(38) => N481, Z(37) => N480, Z(36) => N479, Z(35) => N478, 
               Z(34) => N477, Z(33) => N476, Z(32) => N475, Z(31) => N474, 
               Z(30) => N473, Z(29) => N472, Z(28) => N471, Z(27) => N470, 
               Z(26) => N469, Z(25) => N468, Z(24) => N467, Z(23) => N466, 
               Z(22) => N465, Z(21) => N464, Z(20) => N463, Z(19) => N462, 
               Z(18) => N461, Z(17) => N460, Z(16) => N459, Z(15) => N458, 
               Z(14) => N457, Z(13) => N456, Z(12) => N455, Z(11) => N454, 
               Z(10) => N453, Z(9) => N452, Z(8) => N451, Z(7) => N450, Z(6) =>
               N449, Z(5) => N448, Z(4) => N447, Z(3) => N446, Z(2) => N445, 
               Z(1) => N444, Z(0) => N443 );
   B_28 : GTECH_BUF port map( A => N442, Z => N28);
   B_29 : GTECH_BUF port map( A => state_main_sel(4), Z => N29);
   C1649_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 128 )
      port map(
         -- Connections to port 'DATA1'
         DATA(127) => N570, DATA(126) => N569, DATA(125) => N568, DATA(124) => 
               N567, DATA(123) => N566, DATA(122) => N565, DATA(121) => N564, 
               DATA(120) => N563, DATA(119) => N562, DATA(118) => N561, 
               DATA(117) => N560, DATA(116) => N559, DATA(115) => N558, 
               DATA(114) => N557, DATA(113) => N556, DATA(112) => N555, 
               DATA(111) => N554, DATA(110) => N553, DATA(109) => N552, 
               DATA(108) => N551, DATA(107) => N550, DATA(106) => N549, 
               DATA(105) => N548, DATA(104) => N547, DATA(103) => N546, 
               DATA(102) => N545, DATA(101) => N544, DATA(100) => N543, 
               DATA(99) => N542, DATA(98) => N541, DATA(97) => N540, DATA(96) 
               => N539, DATA(95) => N538, DATA(94) => N537, DATA(93) => N536, 
               DATA(92) => N535, DATA(91) => N534, DATA(90) => N533, DATA(89) 
               => N532, DATA(88) => N531, DATA(87) => N530, DATA(86) => N529, 
               DATA(85) => N528, DATA(84) => N527, DATA(83) => N526, DATA(82) 
               => N525, DATA(81) => N524, DATA(80) => N523, DATA(79) => N522, 
               DATA(78) => N521, DATA(77) => N520, DATA(76) => N519, DATA(75) 
               => N518, DATA(74) => N517, DATA(73) => N516, DATA(72) => N515, 
               DATA(71) => N514, DATA(70) => N513, DATA(69) => N512, DATA(68) 
               => N511, DATA(67) => N510, DATA(66) => N509, DATA(65) => N508, 
               DATA(64) => N507, DATA(63) => N506, DATA(62) => N505, DATA(61) 
               => N504, DATA(60) => N503, DATA(59) => N502, DATA(58) => N501, 
               DATA(57) => N500, DATA(56) => N499, DATA(55) => N498, DATA(54) 
               => N497, DATA(53) => N496, DATA(52) => N495, DATA(51) => N494, 
               DATA(50) => N493, DATA(49) => N492, DATA(48) => N491, DATA(47) 
               => N490, DATA(46) => N489, DATA(45) => N488, DATA(44) => N487, 
               DATA(43) => N486, DATA(42) => N485, DATA(41) => N484, DATA(40) 
               => N483, DATA(39) => N482, DATA(38) => N481, DATA(37) => N480, 
               DATA(36) => N479, DATA(35) => N478, DATA(34) => N477, DATA(33) 
               => N476, DATA(32) => N475, DATA(31) => N474, DATA(30) => N473, 
               DATA(29) => N472, DATA(28) => N471, DATA(27) => N470, DATA(26) 
               => N469, DATA(25) => N468, DATA(24) => N467, DATA(23) => N466, 
               DATA(22) => N465, DATA(21) => N464, DATA(20) => N463, DATA(19) 
               => N462, DATA(18) => N461, DATA(17) => N460, DATA(16) => N459, 
               DATA(15) => N458, DATA(14) => N457, DATA(13) => N456, DATA(12) 
               => N455, DATA(11) => N454, DATA(10) => N453, DATA(9) => N452, 
               DATA(8) => N451, DATA(7) => N450, DATA(6) => N449, DATA(5) => 
               N448, DATA(4) => N447, DATA(3) => N446, DATA(2) => N445, DATA(1)
               => N444, DATA(0) => N443, 
         -- Connections to port 'DATA2'
         DATA(255) => X_Logic0_port, DATA(254) => X_Logic0_port, DATA(253) => 
               X_Logic0_port, DATA(252) => X_Logic0_port, DATA(251) => 
               X_Logic0_port, DATA(250) => X_Logic0_port, DATA(249) => 
               X_Logic0_port, DATA(248) => X_Logic0_port, DATA(247) => 
               X_Logic0_port, DATA(246) => X_Logic0_port, DATA(245) => 
               X_Logic0_port, DATA(244) => X_Logic0_port, DATA(243) => 
               X_Logic0_port, DATA(242) => X_Logic0_port, DATA(241) => 
               X_Logic0_port, DATA(240) => X_Logic0_port, DATA(239) => 
               X_Logic0_port, DATA(238) => X_Logic0_port, DATA(237) => 
               X_Logic0_port, DATA(236) => X_Logic0_port, DATA(235) => 
               X_Logic0_port, DATA(234) => X_Logic0_port, DATA(233) => 
               X_Logic0_port, DATA(232) => X_Logic0_port, DATA(231) => 
               X_Logic0_port, DATA(230) => X_Logic0_port, DATA(229) => 
               X_Logic0_port, DATA(228) => X_Logic0_port, DATA(227) => 
               X_Logic0_port, DATA(226) => X_Logic0_port, DATA(225) => 
               X_Logic0_port, DATA(224) => X_Logic0_port, DATA(223) => 
               X_Logic0_port, DATA(222) => X_Logic0_port, DATA(221) => 
               X_Logic0_port, DATA(220) => X_Logic0_port, DATA(219) => 
               X_Logic0_port, DATA(218) => X_Logic0_port, DATA(217) => 
               X_Logic0_port, DATA(216) => X_Logic0_port, DATA(215) => 
               X_Logic0_port, DATA(214) => X_Logic0_port, DATA(213) => 
               X_Logic0_port, DATA(212) => X_Logic0_port, DATA(211) => 
               X_Logic0_port, DATA(210) => X_Logic0_port, DATA(209) => 
               X_Logic0_port, DATA(208) => X_Logic0_port, DATA(207) => 
               X_Logic0_port, DATA(206) => X_Logic0_port, DATA(205) => 
               X_Logic0_port, DATA(204) => X_Logic0_port, DATA(203) => 
               X_Logic0_port, DATA(202) => X_Logic0_port, DATA(201) => 
               X_Logic0_port, DATA(200) => X_Logic0_port, DATA(199) => 
               X_Logic0_port, DATA(198) => X_Logic0_port, DATA(197) => 
               X_Logic0_port, DATA(196) => X_Logic0_port, DATA(195) => 
               X_Logic0_port, DATA(194) => X_Logic0_port, DATA(193) => 
               X_Logic0_port, DATA(192) => X_Logic0_port, DATA(191) => 
               X_Logic0_port, DATA(190) => X_Logic0_port, DATA(189) => 
               X_Logic0_port, DATA(188) => X_Logic0_port, DATA(187) => 
               X_Logic0_port, DATA(186) => X_Logic0_port, DATA(185) => 
               X_Logic0_port, DATA(184) => X_Logic0_port, DATA(183) => 
               X_Logic0_port, DATA(182) => X_Logic0_port, DATA(181) => 
               X_Logic0_port, DATA(180) => X_Logic0_port, DATA(179) => 
               X_Logic0_port, DATA(178) => X_Logic0_port, DATA(177) => 
               X_Logic0_port, DATA(176) => X_Logic0_port, DATA(175) => 
               X_Logic0_port, DATA(174) => X_Logic0_port, DATA(173) => 
               X_Logic0_port, DATA(172) => X_Logic0_port, DATA(171) => 
               X_Logic0_port, DATA(170) => X_Logic0_port, DATA(169) => 
               X_Logic0_port, DATA(168) => X_Logic0_port, DATA(167) => 
               X_Logic0_port, DATA(166) => X_Logic0_port, DATA(165) => 
               X_Logic0_port, DATA(164) => X_Logic0_port, DATA(163) => 
               X_Logic0_port, DATA(162) => X_Logic0_port, DATA(161) => 
               X_Logic0_port, DATA(160) => X_Logic0_port, DATA(159) => 
               X_Logic0_port, DATA(158) => X_Logic0_port, DATA(157) => 
               X_Logic0_port, DATA(156) => X_Logic0_port, DATA(155) => 
               X_Logic0_port, DATA(154) => X_Logic0_port, DATA(153) => 
               X_Logic0_port, DATA(152) => X_Logic0_port, DATA(151) => 
               X_Logic0_port, DATA(150) => X_Logic0_port, DATA(149) => 
               X_Logic0_port, DATA(148) => X_Logic0_port, DATA(147) => 
               X_Logic0_port, DATA(146) => X_Logic0_port, DATA(145) => 
               X_Logic0_port, DATA(144) => X_Logic0_port, DATA(143) => 
               X_Logic0_port, DATA(142) => X_Logic0_port, DATA(141) => 
               X_Logic0_port, DATA(140) => X_Logic0_port, DATA(139) => 
               X_Logic0_port, DATA(138) => X_Logic0_port, DATA(137) => 
               X_Logic0_port, DATA(136) => X_Logic0_port, DATA(135) => 
               X_Logic0_port, DATA(134) => X_Logic0_port, DATA(133) => 
               X_Logic0_port, DATA(132) => X_Logic0_port, DATA(131) => 
               X_Logic0_port, DATA(130) => X_Logic0_port, DATA(129) => 
               X_Logic0_port, DATA(128) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N30, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N31, 
         -- Connections to port 'Z'
         Z(127) => state_main_in_p2_127_port, Z(126) => 
               state_main_in_p2_126_port, Z(125) => state_main_in_p2_125_port, 
               Z(124) => state_main_in_p2_124_port, Z(123) => 
               state_main_in_p2_123_port, Z(122) => state_main_in_p2_122_port, 
               Z(121) => state_main_in_p2_121_port, Z(120) => 
               state_main_in_p2_120_port, Z(119) => state_main_in_p2_119_port, 
               Z(118) => state_main_in_p2_118_port, Z(117) => 
               state_main_in_p2_117_port, Z(116) => state_main_in_p2_116_port, 
               Z(115) => state_main_in_p2_115_port, Z(114) => 
               state_main_in_p2_114_port, Z(113) => state_main_in_p2_113_port, 
               Z(112) => state_main_in_p2_112_port, Z(111) => 
               state_main_in_p2_111_port, Z(110) => state_main_in_p2_110_port, 
               Z(109) => state_main_in_p2_109_port, Z(108) => 
               state_main_in_p2_108_port, Z(107) => state_main_in_p2_107_port, 
               Z(106) => state_main_in_p2_106_port, Z(105) => 
               state_main_in_p2_105_port, Z(104) => state_main_in_p2_104_port, 
               Z(103) => state_main_in_p2_103_port, Z(102) => 
               state_main_in_p2_102_port, Z(101) => state_main_in_p2_101_port, 
               Z(100) => state_main_in_p2_100_port, Z(99) => 
               state_main_in_p2_99_port, Z(98) => state_main_in_p2_98_port, 
               Z(97) => state_main_in_p2_97_port, Z(96) => 
               state_main_in_p2_96_port, Z(95) => state_main_in_p2_95_port, 
               Z(94) => state_main_in_p2_94_port, Z(93) => 
               state_main_in_p2_93_port, Z(92) => state_main_in_p2_92_port, 
               Z(91) => state_main_in_p2_91_port, Z(90) => 
               state_main_in_p2_90_port, Z(89) => state_main_in_p2_89_port, 
               Z(88) => state_main_in_p2_88_port, Z(87) => 
               state_main_in_p2_87_port, Z(86) => state_main_in_p2_86_port, 
               Z(85) => state_main_in_p2_85_port, Z(84) => 
               state_main_in_p2_84_port, Z(83) => state_main_in_p2_83_port, 
               Z(82) => state_main_in_p2_82_port, Z(81) => 
               state_main_in_p2_81_port, Z(80) => state_main_in_p2_80_port, 
               Z(79) => state_main_in_p2_79_port, Z(78) => 
               state_main_in_p2_78_port, Z(77) => state_main_in_p2_77_port, 
               Z(76) => state_main_in_p2_76_port, Z(75) => 
               state_main_in_p2_75_port, Z(74) => state_main_in_p2_74_port, 
               Z(73) => state_main_in_p2_73_port, Z(72) => 
               state_main_in_p2_72_port, Z(71) => state_main_in_p2_71_port, 
               Z(70) => state_main_in_p2_70_port, Z(69) => 
               state_main_in_p2_69_port, Z(68) => state_main_in_p2_68_port, 
               Z(67) => state_main_in_p2_67_port, Z(66) => 
               state_main_in_p2_66_port, Z(65) => state_main_in_p2_65_port, 
               Z(64) => state_main_in_p2_64_port, Z(63) => 
               state_main_in_p2_63_port, Z(62) => state_main_in_p2_62_port, 
               Z(61) => state_main_in_p2_61_port, Z(60) => 
               state_main_in_p2_60_port, Z(59) => state_main_in_p2_59_port, 
               Z(58) => state_main_in_p2_58_port, Z(57) => 
               state_main_in_p2_57_port, Z(56) => state_main_in_p2_56_port, 
               Z(55) => state_main_in_p2_55_port, Z(54) => 
               state_main_in_p2_54_port, Z(53) => state_main_in_p2_53_port, 
               Z(52) => state_main_in_p2_52_port, Z(51) => 
               state_main_in_p2_51_port, Z(50) => state_main_in_p2_50_port, 
               Z(49) => state_main_in_p2_49_port, Z(48) => 
               state_main_in_p2_48_port, Z(47) => state_main_in_p2_47_port, 
               Z(46) => state_main_in_p2_46_port, Z(45) => 
               state_main_in_p2_45_port, Z(44) => state_main_in_p2_44_port, 
               Z(43) => state_main_in_p2_43_port, Z(42) => 
               state_main_in_p2_42_port, Z(41) => state_main_in_p2_41_port, 
               Z(40) => state_main_in_p2_40_port, Z(39) => 
               state_main_in_p2_39_port, Z(38) => state_main_in_p2_38_port, 
               Z(37) => state_main_in_p2_37_port, Z(36) => 
               state_main_in_p2_36_port, Z(35) => state_main_in_p2_35_port, 
               Z(34) => state_main_in_p2_34_port, Z(33) => 
               state_main_in_p2_33_port, Z(32) => state_main_in_p2_32_port, 
               Z(31) => state_main_in_p2_31_port, Z(30) => 
               state_main_in_p2_30_port, Z(29) => state_main_in_p2_29_port, 
               Z(28) => state_main_in_p2_28_port, Z(27) => 
               state_main_in_p2_27_port, Z(26) => state_main_in_p2_26_port, 
               Z(25) => state_main_in_p2_25_port, Z(24) => 
               state_main_in_p2_24_port, Z(23) => state_main_in_p2_23_port, 
               Z(22) => state_main_in_p2_22_port, Z(21) => 
               state_main_in_p2_21_port, Z(20) => state_main_in_p2_20_port, 
               Z(19) => state_main_in_p2_19_port, Z(18) => 
               state_main_in_p2_18_port, Z(17) => state_main_in_p2_17_port, 
               Z(16) => state_main_in_p2_16_port, Z(15) => 
               state_main_in_p2_15_port, Z(14) => state_main_in_p2_14_port, 
               Z(13) => state_main_in_p2_13_port, Z(12) => 
               state_main_in_p2_12_port, Z(11) => state_main_in_p2_11_port, 
               Z(10) => state_main_in_p2_10_port, Z(9) => 
               state_main_in_p2_9_port, Z(8) => state_main_in_p2_8_port, Z(7) 
               => state_main_in_p2_7_port, Z(6) => state_main_in_p2_6_port, 
               Z(5) => state_main_in_p2_5_port, Z(4) => state_main_in_p2_4_port
               , Z(3) => state_main_in_p2_3_port, Z(2) => 
               state_main_in_p2_2_port, Z(1) => state_main_in_p2_1_port, Z(0) 
               => state_main_in_p2_0_port );
   B_30 : GTECH_BUF port map( A => N441, Z => N30);
   B_31 : GTECH_BUF port map( A => state_main_sel(5), Z => N31);
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   I_4 : GTECH_NOT port map( A => dcount_in(3), Z => N32);
   I_5 : GTECH_NOT port map( A => dcount_in(2), Z => N33);
   I_6 : GTECH_NOT port map( A => N162, Z => N163);
   I_7 : GTECH_NOT port map( A => N164, Z => N165);
   I_8 : GTECH_NOT port map( A => cycd_sel(1), Z => N167);
   I_9 : GTECH_NOT port map( A => cycd_sel(0), Z => N168);
   C1668 : GTECH_XOR2 port map( A => temp_ram_31_port, B => xor_mux_o_31_port, 
                           Z => temp_xor_out_31_port);
   C1669 : GTECH_XOR2 port map( A => temp_ram_30_port, B => xor_mux_o_30_port, 
                           Z => temp_xor_out_30_port);
   C1670 : GTECH_XOR2 port map( A => temp_ram_29_port, B => xor_mux_o_29_port, 
                           Z => temp_xor_out_29_port);
   C1671 : GTECH_XOR2 port map( A => temp_ram_28_port, B => xor_mux_o_28_port, 
                           Z => temp_xor_out_28_port);
   C1672 : GTECH_XOR2 port map( A => temp_ram_27_port, B => xor_mux_o_27_port, 
                           Z => temp_xor_out_27_port);
   C1673 : GTECH_XOR2 port map( A => temp_ram_26_port, B => xor_mux_o_26_port, 
                           Z => temp_xor_out_26_port);
   C1674 : GTECH_XOR2 port map( A => temp_ram_25_port, B => xor_mux_o_25_port, 
                           Z => temp_xor_out_25_port);
   C1675 : GTECH_XOR2 port map( A => temp_ram_24_port, B => xor_mux_o_24_port, 
                           Z => temp_xor_out_24_port);
   C1676 : GTECH_XOR2 port map( A => temp_ram_23_port, B => xor_mux_o_23_port, 
                           Z => temp_xor_out_23_port);
   C1677 : GTECH_XOR2 port map( A => temp_ram_22_port, B => xor_mux_o_22_port, 
                           Z => temp_xor_out_22_port);
   C1678 : GTECH_XOR2 port map( A => temp_ram_21_port, B => xor_mux_o_21_port, 
                           Z => temp_xor_out_21_port);
   C1679 : GTECH_XOR2 port map( A => temp_ram_20_port, B => xor_mux_o_20_port, 
                           Z => temp_xor_out_20_port);
   C1680 : GTECH_XOR2 port map( A => temp_ram_19_port, B => xor_mux_o_19_port, 
                           Z => temp_xor_out_19_port);
   C1681 : GTECH_XOR2 port map( A => temp_ram_18_port, B => xor_mux_o_18_port, 
                           Z => temp_xor_out_18_port);
   C1682 : GTECH_XOR2 port map( A => temp_ram_17_port, B => xor_mux_o_17_port, 
                           Z => temp_xor_out_17_port);
   C1683 : GTECH_XOR2 port map( A => temp_ram_16_port, B => xor_mux_o_16_port, 
                           Z => temp_xor_out_16_port);
   C1684 : GTECH_XOR2 port map( A => temp_ram_15_port, B => xor_mux_o_15_port, 
                           Z => temp_xor_out_15_port);
   C1685 : GTECH_XOR2 port map( A => temp_ram_14_port, B => xor_mux_o_14_port, 
                           Z => temp_xor_out_14_port);
   C1686 : GTECH_XOR2 port map( A => temp_ram_13_port, B => xor_mux_o_13_port, 
                           Z => temp_xor_out_13_port);
   C1687 : GTECH_XOR2 port map( A => temp_ram_12_port, B => xor_mux_o_12_port, 
                           Z => temp_xor_out_12_port);
   C1688 : GTECH_XOR2 port map( A => temp_ram_11_port, B => xor_mux_o_11_port, 
                           Z => temp_xor_out_11_port);
   C1689 : GTECH_XOR2 port map( A => temp_ram_10_port, B => xor_mux_o_10_port, 
                           Z => temp_xor_out_10_port);
   C1690 : GTECH_XOR2 port map( A => temp_ram_9_port, B => xor_mux_o_9_port, Z 
                           => temp_xor_out_9_port);
   C1691 : GTECH_XOR2 port map( A => temp_ram_8_port, B => xor_mux_o_8_port, Z 
                           => temp_xor_out_8_port);
   C1692 : GTECH_XOR2 port map( A => temp_ram_7_port, B => xor_mux_o_7_port, Z 
                           => temp_xor_out_7_port);
   C1693 : GTECH_XOR2 port map( A => temp_ram_6_port, B => xor_mux_o_6_port, Z 
                           => temp_xor_out_6_port);
   C1694 : GTECH_XOR2 port map( A => temp_ram_5_port, B => xor_mux_o_5_port, Z 
                           => temp_xor_out_5_port);
   C1695 : GTECH_XOR2 port map( A => temp_ram_4_port, B => xor_mux_o_4_port, Z 
                           => temp_xor_out_4_port);
   C1696 : GTECH_XOR2 port map( A => temp_ram_3_port, B => xor_mux_o_3_port, Z 
                           => temp_xor_out_3_port);
   C1697 : GTECH_XOR2 port map( A => temp_ram_2_port, B => xor_mux_o_2_port, Z 
                           => temp_xor_out_2_port);
   C1698 : GTECH_XOR2 port map( A => temp_ram_1_port, B => xor_mux_o_1_port, Z 
                           => temp_xor_out_1_port);
   C1699 : GTECH_XOR2 port map( A => temp_ram_0_port, B => xor_mux_o_0_port, Z 
                           => temp_xor_out_0_port);
   I_10 : GTECH_NOT port map( A => dcount_in(1), Z => N170);
   I_11 : GTECH_NOT port map( A => dcount_in(0), Z => N171);
   I_12 : GTECH_NOT port map( A => N173, Z => N174);
   I_13 : GTECH_NOT port map( A => N175, Z => N176);
   I_14 : GTECH_NOT port map( A => temp_ram_8_port, Z => N178);
   I_15 : GTECH_NOT port map( A => temp_ram_16_port, Z => N179);
   I_16 : GTECH_NOT port map( A => temp_ram_24_port, Z => N180);
   C1719 : GTECH_XOR2 port map( A => state_main_out_plane2_31_port, B => 
                           cu_cd(7), Z => fb_prime_7_port);
   C1720 : GTECH_XOR2 port map( A => state_main_out_plane2_30_port, B => 
                           cu_cd(6), Z => fb_prime_6_port);
   C1721 : GTECH_XOR2 port map( A => state_main_out_plane2_29_port, B => 
                           cu_cd(5), Z => fb_prime_5_port);
   C1722 : GTECH_XOR2 port map( A => state_main_out_plane2_28_port, B => 
                           cu_cd(4), Z => fb_prime_4_port);
   C1723 : GTECH_XOR2 port map( A => state_main_out_plane2_27_port, B => 
                           cu_cd(3), Z => fb_prime_3_port);
   C1724 : GTECH_XOR2 port map( A => state_main_out_plane2_26_port, B => 
                           cu_cd(2), Z => fb_prime_2_port);
   C1725 : GTECH_XOR2 port map( A => state_main_out_plane2_25_port, B => 
                           cu_cd(1), Z => fb_prime_1_port);
   C1726 : GTECH_XOR2 port map( A => state_main_out_plane2_24_port, B => 
                           cu_cd(0), Z => fb_prime_0_port);
   I_17 : GTECH_NOT port map( A => state_main_sel(1), Z => N181);
   I_18 : GTECH_NOT port map( A => state_main_sel(0), Z => N182);
   I_19 : GTECH_NOT port map( A => state_main_sel(3), Z => N311);
   I_20 : GTECH_NOT port map( A => state_main_sel(2), Z => N312);
   I_21 : GTECH_NOT port map( A => state_main_sel(5), Z => N441);
   I_22 : GTECH_NOT port map( A => state_main_sel(4), Z => N442);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_LWC_1.all;

entity counter_num_bits4_1 is

   port( clk, reset, enable : in std_logic;  q : out std_logic_vector (3 downto
         0));

end counter_num_bits4_1;

architecture SYN_Behavioral of counter_num_bits4_1 is

   component GTECH_AND2
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component GTECH_BUF
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component GTECH_NOT
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
      generic ( ac_as_q, ac_as_qn, sc_ss_q : integer );
      port(
         clear, preset, enable, data_in, synch_clear, synch_preset, 
            synch_toggle, synch_enable, next_state, clocked_on : in std_logic;
         Q, QN : buffer std_logic
      );
   end component;
   
   signal N0, N1, X_Logic1_port, X_Logic0_port, clk_port, enable_port, q_3_port
      , q_2_port, q_1_port, q_0_port, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11,
      N12, n_1128, n_1129, n_1130, n_1131, n_1132 : std_logic;

begin
   clk_port <= clk;
   enable_port <= enable;
   q <= ( q_3_port, q_2_port, q_1_port, q_0_port );
   
   count_reg_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N8, next_state => N12, clocked_on
               => clk_port, Q => q_3_port, QN => n_1128);
   count_reg_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N8, next_state => N11, clocked_on
               => clk_port, Q => q_2_port, QN => n_1129);
   count_reg_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N8, next_state => N10, clocked_on
               => clk_port, Q => q_1_port, QN => n_1130);
   count_reg_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N8, next_state => N9, clocked_on 
               => clk_port, Q => q_0_port, QN => n_1131);
   add_39 : process ( q_3_port, q_2_port, q_1_port, q_0_port, X_Logic1_port )
      variable A : UNSIGNED( 3 downto 0 );
      variable B : UNSIGNED( 3 downto 0 );
      variable Z : UNSIGNED( 3 downto 0 );
   begin
      A := ( q_3_port, q_2_port, q_1_port, q_0_port );
      B := ( '0', '0', '0', X_Logic1_port );
      Z := A + B;
      ( N7, N6, N5, N4 ) <= Z;
   end process;
   
   C33_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic1_port, 
         -- Connections to port 'DATA2'
         DATA(1) => enable_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N0, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N1, 
         -- Connections to port 'Z'
         Z(0) => N8 );
   B_0 : GTECH_BUF port map( A => reset, Z => N0);
   B_1 : GTECH_BUF port map( A => N2, Z => N1);
   C34_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 4 )
      port map(
         -- Connections to port 'DATA1'
         DATA(3) => X_Logic0_port, DATA(2) => X_Logic0_port, DATA(1) => 
               X_Logic0_port, DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(7) => N7, DATA(6) => N6, DATA(5) => N5, DATA(4) => N4, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N0, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N1, 
         -- Connections to port 'Z'
         Z(3) => N12, Z(2) => N11, Z(1) => N10, Z(0) => N9 );
         X_Logic1_port <= '1';
         X_Logic0_port <= '0';
   I_0 : GTECH_NOT port map( A => reset, Z => N2);
   B_2 : GTECH_BUF port map( A => N2, Z => N3);
   C42 : GTECH_AND2 port map( A => N3, B => enable_port, Z => n_1132);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_LWC_1.all;

entity DATA_PISO_2 is

   port( clk, rst : in std_logic;  data_size_p : in std_logic_vector (2 downto 
         0);  data_size_s : out std_logic_vector (2 downto 0);  data_s : out 
         std_logic_vector (31 downto 0);  data_valid_s : out std_logic;  
         data_ready_s : in std_logic;  data_p : in std_logic_vector (31 downto 
         0);  data_valid_p : in std_logic;  data_ready_p : out std_logic;  
         valid_bytes_p : in std_logic_vector (3 downto 0);  valid_bytes_s : out
         std_logic_vector (3 downto 0);  pad_loc_p : in std_logic_vector (3 
         downto 0);  pad_loc_s : out std_logic_vector (3 downto 0);  eoi_p : in
         std_logic;  eoi_s : out std_logic;  eot_p : in std_logic;  eot_s : out
         std_logic);

end DATA_PISO_2;

architecture SYN_behavioral of DATA_PISO_2 is

begin
   data_size_s <= ( data_size_p(2), data_size_p(1), data_size_p(0) );
   data_s <= ( data_p(31), data_p(30), data_p(29), data_p(28), data_p(27), 
      data_p(26), data_p(25), data_p(24), data_p(23), data_p(22), data_p(21), 
      data_p(20), data_p(19), data_p(18), data_p(17), data_p(16), data_p(15), 
      data_p(14), data_p(13), data_p(12), data_p(11), data_p(10), data_p(9), 
      data_p(8), data_p(7), data_p(6), data_p(5), data_p(4), data_p(3), 
      data_p(2), data_p(1), data_p(0) );
   data_valid_s <= data_valid_p;
   data_ready_p <= data_ready_s;
   valid_bytes_s <= ( valid_bytes_p(3), valid_bytes_p(2), valid_bytes_p(1), 
      valid_bytes_p(0) );
   pad_loc_s <= ( pad_loc_p(3), pad_loc_p(2), pad_loc_p(1), pad_loc_p(0) );
   eoi_s <= eoi_p;
   eot_s <= eot_p;

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_LWC_1.all;

entity KEY_PISO_2 is

   port( clk, rst : in std_logic;  data_s : out std_logic_vector (31 downto 0);
         data_valid_s : out std_logic;  data_ready_s : in std_logic;  data_p : 
         in std_logic_vector (31 downto 0);  data_valid_p : in std_logic;  
         data_ready_p : out std_logic);

end KEY_PISO_2;

architecture SYN_behavioral of KEY_PISO_2 is

begin
   data_s <= ( data_p(31), data_p(30), data_p(29), data_p(28), data_p(27), 
      data_p(26), data_p(25), data_p(24), data_p(23), data_p(22), data_p(21), 
      data_p(20), data_p(19), data_p(18), data_p(17), data_p(16), data_p(15), 
      data_p(14), data_p(13), data_p(12), data_p(11), data_p(10), data_p(9), 
      data_p(8), data_p(7), data_p(6), data_p(5), data_p(4), data_p(3), 
      data_p(2), data_p(1), data_p(0) );
   data_valid_s <= data_valid_p;
   data_ready_p <= data_ready_s;

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_LWC_1.all;

entity StepDownCountLd_N16_step4_2 is

   port( clk, len, ena : in std_logic;  load : in std_logic_vector (15 downto 
         0);  count : out std_logic_vector (15 downto 0));

end StepDownCountLd_N16_step4_2;

architecture SYN_StepDownCountLd of StepDownCountLd_N16_step4_2 is

   component GTECH_AND2
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component GTECH_BUF
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component GTECH_NOT
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
      generic ( ac_as_q, ac_as_qn, sc_ss_q : integer );
      port(
         clear, preset, enable, data_in, synch_clear, synch_preset, 
            synch_toggle, synch_enable, next_state, clocked_on : in std_logic;
         Q, QN : buffer std_logic
      );
   end component;
   
   signal N0, N1, X_Logic1_port, X_Logic0_port, clk_port, ena_port, 
      load_15_port, load_14_port, load_13_port, load_12_port, load_11_port, 
      load_10_port, load_9_port, load_8_port, load_7_port, load_6_port, 
      load_5_port, load_4_port, load_3_port, load_2_port, load_1_port, 
      load_0_port, count_15_port, count_14_port, count_13_port, count_12_port, 
      count_11_port, count_10_port, count_9_port, count_8_port, count_7_port, 
      count_6_port, count_5_port, count_4_port, count_3_port, count_2_port, 
      count_1_port, count_0_port, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12
      , N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, 
      N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, n_1133, n_1134, n_1135,
      n_1136, n_1137, n_1138, n_1139, n_1140, n_1141, n_1142, n_1143, n_1144, 
      n_1145, n_1146, n_1147, n_1148, n_1149 : std_logic;

begin
   clk_port <= clk;
   ena_port <= ena;
   ( load_15_port, load_14_port, load_13_port, load_12_port, load_11_port, 
      load_10_port, load_9_port, load_8_port, load_7_port, load_6_port, 
      load_5_port, load_4_port, load_3_port, load_2_port, load_1_port, 
      load_0_port ) <= load;
   count <= ( count_15_port, count_14_port, count_13_port, count_12_port, 
      count_11_port, count_10_port, count_9_port, count_8_port, count_7_port, 
      count_6_port, count_5_port, count_4_port, count_3_port, count_2_port, 
      count_1_port, count_0_port );
   
   qtemp_reg_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N20, next_state => N36, 
               clocked_on => clk_port, Q => count_15_port, QN => n_1133);
   qtemp_reg_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N20, next_state => N35, 
               clocked_on => clk_port, Q => count_14_port, QN => n_1134);
   qtemp_reg_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N20, next_state => N34, 
               clocked_on => clk_port, Q => count_13_port, QN => n_1135);
   qtemp_reg_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N20, next_state => N33, 
               clocked_on => clk_port, Q => count_12_port, QN => n_1136);
   qtemp_reg_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N20, next_state => N32, 
               clocked_on => clk_port, Q => count_11_port, QN => n_1137);
   qtemp_reg_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N20, next_state => N31, 
               clocked_on => clk_port, Q => count_10_port, QN => n_1138);
   qtemp_reg_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N20, next_state => N30, 
               clocked_on => clk_port, Q => count_9_port, QN => n_1139);
   qtemp_reg_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N20, next_state => N29, 
               clocked_on => clk_port, Q => count_8_port, QN => n_1140);
   qtemp_reg_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N20, next_state => N28, 
               clocked_on => clk_port, Q => count_7_port, QN => n_1141);
   qtemp_reg_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N20, next_state => N27, 
               clocked_on => clk_port, Q => count_6_port, QN => n_1142);
   qtemp_reg_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N20, next_state => N26, 
               clocked_on => clk_port, Q => count_5_port, QN => n_1143);
   qtemp_reg_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N20, next_state => N25, 
               clocked_on => clk_port, Q => count_4_port, QN => n_1144);
   qtemp_reg_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N20, next_state => N24, 
               clocked_on => clk_port, Q => count_3_port, QN => n_1145);
   qtemp_reg_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N20, next_state => N23, 
               clocked_on => clk_port, Q => count_2_port, QN => n_1146);
   qtemp_reg_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N20, next_state => N22, 
               clocked_on => clk_port, Q => count_1_port, QN => n_1147);
   qtemp_reg_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N20, next_state => N21, 
               clocked_on => clk_port, Q => count_0_port, QN => n_1148);
   sub_55 : process ( count_15_port, count_14_port, count_13_port, 
         count_12_port, count_11_port, count_10_port, count_9_port, 
         count_8_port, count_7_port, count_6_port, count_5_port, count_4_port, 
         count_3_port, count_2_port, count_1_port, count_0_port, X_Logic1_port,
         X_Logic0_port )
      variable A : UNSIGNED( 15 downto 0 );
      variable B : UNSIGNED( 15 downto 0 );
      variable Z : UNSIGNED( 15 downto 0 );
   begin
      A := ( count_15_port, count_14_port, count_13_port, count_12_port, 
            count_11_port, count_10_port, count_9_port, count_8_port, 
            count_7_port, count_6_port, count_5_port, count_4_port, 
            count_3_port, count_2_port, count_1_port, count_0_port );
      B := ( '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', 
            X_Logic1_port, X_Logic0_port, X_Logic0_port );
      Z := A - B;
      ( N19, N18, N17, N16, N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, 
            N4 ) <= Z;
   end process;
   
   C81_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic1_port, 
         -- Connections to port 'DATA2'
         DATA(1) => ena_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N0, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N1, 
         -- Connections to port 'Z'
         Z(0) => N20 );
   B_0 : GTECH_BUF port map( A => len, Z => N0);
   B_1 : GTECH_BUF port map( A => N2, Z => N1);
   C82_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 16 )
      port map(
         -- Connections to port 'DATA1'
         DATA(15) => load_15_port, DATA(14) => load_14_port, DATA(13) => 
               load_13_port, DATA(12) => load_12_port, DATA(11) => load_11_port
               , DATA(10) => load_10_port, DATA(9) => load_9_port, DATA(8) => 
               load_8_port, DATA(7) => load_7_port, DATA(6) => load_6_port, 
               DATA(5) => load_5_port, DATA(4) => load_4_port, DATA(3) => 
               load_3_port, DATA(2) => load_2_port, DATA(1) => load_1_port, 
               DATA(0) => load_0_port, 
         -- Connections to port 'DATA2'
         DATA(31) => N19, DATA(30) => N18, DATA(29) => N17, DATA(28) => N16, 
               DATA(27) => N15, DATA(26) => N14, DATA(25) => N13, DATA(24) => 
               N12, DATA(23) => N11, DATA(22) => N10, DATA(21) => N9, DATA(20) 
               => N8, DATA(19) => N7, DATA(18) => N6, DATA(17) => N5, DATA(16) 
               => N4, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N0, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N1, 
         -- Connections to port 'Z'
         Z(15) => N36, Z(14) => N35, Z(13) => N34, Z(12) => N33, Z(11) => N32, 
               Z(10) => N31, Z(9) => N30, Z(8) => N29, Z(7) => N28, Z(6) => N27
               , Z(5) => N26, Z(4) => N25, Z(3) => N24, Z(2) => N23, Z(1) => 
               N22, Z(0) => N21 );
         X_Logic1_port <= '1';
         X_Logic0_port <= '0';
   I_0 : GTECH_NOT port map( A => len, Z => N2);
   B_2 : GTECH_BUF port map( A => N2, Z => N3);
   C90 : GTECH_AND2 port map( A => N3, B => ena_port, Z => n_1149);

end SYN_StepDownCountLd;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_LWC_1.all;

entity PostProcessor_2 is

   port( clk, rst : in std_logic;  bdo : in std_logic_vector (31 downto 0);  
         bdo_valid : in std_logic;  bdo_ready : out std_logic;  end_of_block : 
         in std_logic;  bdo_type, bdo_valid_bytes : in std_logic_vector (3 
         downto 0);  msg_auth : in std_logic;  msg_auth_ready : out std_logic; 
         msg_auth_valid : in std_logic;  cmd : in std_logic_vector (31 downto 
         0);  cmd_valid : in std_logic;  cmd_ready : out std_logic;  do_data : 
         out std_logic_vector (31 downto 0);  do_valid, do_last : out std_logic
         ;  do_ready : in std_logic);

end PostProcessor_2;

architecture SYN_PostProcessor of PostProcessor_2 is

   component GTECH_NOT
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component GTECH_AND2
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component GTECH_OR2
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component GTECH_BUF
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
      generic ( ac_as_q, ac_as_qn, sc_ss_q : integer );
      port(
         clear, preset, enable, data_in, synch_clear, synch_preset, 
            synch_toggle, synch_enable, next_state, clocked_on : in std_logic;
         Q, QN : buffer std_logic
      );
   end component;
   
   component DATA_SIPO_2
      port( clk, rst, end_of_input : in std_logic;  data_p : out 
            std_logic_vector (31 downto 0);  data_valid_p : out std_logic;  
            data_ready_p : in std_logic;  data_s : in std_logic_vector (31 
            downto 0);  data_valid_s : in std_logic;  data_ready_s : out 
            std_logic);
   end component;
   
   component StepDownCountLd_N16_step4_2
      port( clk, len, ena : in std_logic;  load : in std_logic_vector (15 
            downto 0);  count : out std_logic_vector (15 downto 0));
   end component;
   
   signal N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15,
      N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30
      , N31, N32, N33, N34, N35, N36, N37, N38, X_Logic1_port, X_Logic0_port, 
      clk_port, msg_auth_port, msg_auth_ready_port, msg_auth_valid_port, cmd_31
      , cmd_30, cmd_29, cmd_28, cmd_25, cmd_15_port, cmd_14_port, cmd_13_port, 
      cmd_12_port, cmd_11_port, cmd_10_port, cmd_9_port, cmd_8_port, cmd_7_port
      , cmd_6_port, cmd_5_port, cmd_4_port, cmd_3_port, cmd_2_port, cmd_1_port,
      cmd_0_port, cmd_valid_port, cmd_ready_port, do_data_31_port, 
      do_data_30_port, do_data_29_port, do_data_28_port, do_data_27_port, 
      do_data_26_port, do_data_25_port, do_data_24_port, do_data_23_port, 
      do_data_22_port, do_data_21_port, do_data_20_port, do_data_19_port, 
      do_data_18_port, do_data_17_port, do_data_16_port, do_data_15_port, 
      do_data_14_port, do_data_13_port, do_data_12_port, do_data_11_port, 
      do_data_10_port, do_data_9_port, do_data_8_port, do_data_7_port, 
      do_data_6_port, do_data_5_port, do_data_4_port, do_data_3_port, 
      do_data_2_port, do_data_1_port, do_data_0_port, do_valid_port, 
      do_last_port, do_ready_port, bdo_cleared_31_port, bdo_cleared_30_port, 
      bdo_cleared_29_port, bdo_cleared_28_port, bdo_cleared_27_port, 
      bdo_cleared_26_port, bdo_cleared_25_port, bdo_cleared_24_port, 
      bdo_cleared_23_port, bdo_cleared_22_port, bdo_cleared_21_port, 
      bdo_cleared_20_port, bdo_cleared_19_port, bdo_cleared_18_port, 
      bdo_cleared_17_port, bdo_cleared_16_port, bdo_cleared_15_port, 
      bdo_cleared_14_port, bdo_cleared_13_port, bdo_cleared_12_port, 
      bdo_cleared_11_port, bdo_cleared_10_port, bdo_cleared_9_port, 
      bdo_cleared_8_port, bdo_cleared_7_port, bdo_cleared_6_port, 
      bdo_cleared_5_port, bdo_cleared_4_port, bdo_cleared_3_port, 
      bdo_cleared_2_port, bdo_cleared_1_port, bdo_cleared_0_port, N39, 
      do_data_internal_31_port, do_data_internal_30_port, 
      do_data_internal_29_port, do_data_internal_28_port, 
      do_data_internal_27_port, do_data_internal_26_port, 
      do_data_internal_25_port, do_data_internal_24_port, 
      do_data_internal_23_port, do_data_internal_22_port, 
      do_data_internal_21_port, do_data_internal_20_port, 
      do_data_internal_19_port, do_data_internal_18_port, 
      do_data_internal_17_port, do_data_internal_16_port, 
      do_data_internal_15_port, do_data_internal_14_port, 
      do_data_internal_13_port, do_data_internal_12_port, 
      do_data_internal_11_port, do_data_internal_10_port, 
      do_data_internal_9_port, do_data_internal_8_port, do_data_internal_7_port
      , do_data_internal_6_port, do_data_internal_5_port, 
      do_data_internal_4_port, do_data_internal_3_port, do_data_internal_2_port
      , do_data_internal_1_port, do_data_internal_0_port, len_SegLenCnt, 
      en_SegLenCnt, dout_SegLenCnt_15_port, dout_SegLenCnt_14_port, 
      dout_SegLenCnt_13_port, dout_SegLenCnt_12_port, dout_SegLenCnt_11_port, 
      dout_SegLenCnt_10_port, dout_SegLenCnt_9_port, dout_SegLenCnt_8_port, 
      dout_SegLenCnt_7_port, dout_SegLenCnt_6_port, dout_SegLenCnt_5_port, 
      dout_SegLenCnt_4_port, dout_SegLenCnt_3_port, dout_SegLenCnt_2_port, 
      dout_SegLenCnt_1_port, dout_SegLenCnt_0_port, N40, last_flit_of_segment, 
      eot, decrypt, bdo_ready_p, bdo_valid_p, bdo_p_31_port, bdo_p_30_port, 
      bdo_p_29_port, bdo_p_28_port, bdo_p_27_port, bdo_p_26_port, bdo_p_25_port
      , bdo_p_24_port, bdo_p_23_port, bdo_p_22_port, bdo_p_21_port, 
      bdo_p_20_port, bdo_p_19_port, bdo_p_18_port, bdo_p_17_port, bdo_p_16_port
      , bdo_p_15_port, bdo_p_14_port, bdo_p_13_port, bdo_p_12_port, 
      bdo_p_11_port, bdo_p_10_port, bdo_p_9_port, bdo_p_8_port, bdo_p_7_port, 
      bdo_p_6_port, bdo_p_5_port, bdo_p_4_port, bdo_p_3_port, bdo_p_2_port, 
      bdo_p_1_port, bdo_p_0_port, N41, pr_state_3_port, pr_state_2_port, 
      pr_state_1_port, pr_state_0_port, nx_state_3_port, nx_state_2_port, 
      nx_state_1_port, nx_state_0_port, N42, N43, N44, N45, N46, N47, N48, N49,
      N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64
      , N65, N66, N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78, 
      N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91, N92, N93
      , N94, N95, N96, N97, N98, N99, N100, N101, N102, N103, N104, N105, N106,
      N107, N108, N109, N110, N111, N112, N113, N114, N115, N116, N117, N118, 
      N119, N120, N121, N122, N123, N124, N125, N126, N127, N128, N129, N130, 
      N131, N132, N133, N134, N135, N136, N137, N138, N139, N140, N141, N142, 
      N143, N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154, 
      N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165, N166, 
      N167, N168, N169, N170, N171, N172, N173, N174, N175, N176, N177, N178, 
      N179, N180, N181, N182, N183, N184, N185, N186, N187, N188, N189, N190, 
      N191, N192, N193, N194, N195, N196, N197, N198, N199, N200, N201, N202, 
      N203, N204, N205, N206, net1438, net1439, net1440, net1441, net1442, 
      net1443, net1444, net1445, net1446, net1447, net1448, n_1150, n_1151, 
      n_1152, n_1153, n_1154, n_1155 : std_logic;

begin
   clk_port <= clk;
   msg_auth_port <= msg_auth;
   msg_auth_ready <= msg_auth_ready_port;
   msg_auth_valid_port <= msg_auth_valid;
   ( cmd_31, cmd_30, cmd_29, cmd_28, net1438, net1439, cmd_25, net1440, net1441
      , net1442, net1443, net1444, net1445, net1446, net1447, net1448, 
      cmd_15_port, cmd_14_port, cmd_13_port, cmd_12_port, cmd_11_port, 
      cmd_10_port, cmd_9_port, cmd_8_port, cmd_7_port, cmd_6_port, cmd_5_port, 
      cmd_4_port, cmd_3_port, cmd_2_port, cmd_1_port, cmd_0_port ) <= cmd;
   cmd_valid_port <= cmd_valid;
   cmd_ready <= cmd_ready_port;
   do_data <= ( do_data_31_port, do_data_30_port, do_data_29_port, 
      do_data_28_port, do_data_27_port, do_data_26_port, do_data_25_port, 
      do_data_24_port, do_data_23_port, do_data_22_port, do_data_21_port, 
      do_data_20_port, do_data_19_port, do_data_18_port, do_data_17_port, 
      do_data_16_port, do_data_15_port, do_data_14_port, do_data_13_port, 
      do_data_12_port, do_data_11_port, do_data_10_port, do_data_9_port, 
      do_data_8_port, do_data_7_port, do_data_6_port, do_data_5_port, 
      do_data_4_port, do_data_3_port, do_data_2_port, do_data_1_port, 
      do_data_0_port );
   do_valid <= do_valid_port;
   do_last <= do_last_port;
   do_ready_port <= do_ready;
   
   SegLen : StepDownCountLd_N16_step4_2 port map( clk => clk_port, len => 
                           len_SegLenCnt, ena => en_SegLenCnt, load(15) => 
                           cmd_15_port, load(14) => cmd_14_port, load(13) => 
                           cmd_13_port, load(12) => cmd_12_port, load(11) => 
                           cmd_11_port, load(10) => cmd_10_port, load(9) => 
                           cmd_9_port, load(8) => cmd_8_port, load(7) => 
                           cmd_7_port, load(6) => cmd_6_port, load(5) => 
                           cmd_5_port, load(4) => cmd_4_port, load(3) => 
                           cmd_3_port, load(2) => cmd_2_port, load(1) => 
                           cmd_1_port, load(0) => cmd_0_port, count(15) => 
                           dout_SegLenCnt_15_port, count(14) => 
                           dout_SegLenCnt_14_port, count(13) => 
                           dout_SegLenCnt_13_port, count(12) => 
                           dout_SegLenCnt_12_port, count(11) => 
                           dout_SegLenCnt_11_port, count(10) => 
                           dout_SegLenCnt_10_port, count(9) => 
                           dout_SegLenCnt_9_port, count(8) => 
                           dout_SegLenCnt_8_port, count(7) => 
                           dout_SegLenCnt_7_port, count(6) => 
                           dout_SegLenCnt_6_port, count(5) => 
                           dout_SegLenCnt_5_port, count(4) => 
                           dout_SegLenCnt_4_port, count(3) => 
                           dout_SegLenCnt_3_port, count(2) => 
                           dout_SegLenCnt_2_port, count(1) => 
                           dout_SegLenCnt_1_port, count(0) => 
                           dout_SegLenCnt_0_port);
   lte_146 : process ( dout_SegLenCnt_15_port, dout_SegLenCnt_14_port, 
         dout_SegLenCnt_13_port, dout_SegLenCnt_12_port, dout_SegLenCnt_11_port
         , dout_SegLenCnt_10_port, dout_SegLenCnt_9_port, dout_SegLenCnt_8_port
         , dout_SegLenCnt_7_port, dout_SegLenCnt_6_port, dout_SegLenCnt_5_port,
         dout_SegLenCnt_4_port, dout_SegLenCnt_3_port, dout_SegLenCnt_2_port, 
         dout_SegLenCnt_1_port, dout_SegLenCnt_0_port, X_Logic0_port, 
         X_Logic1_port )
      variable A : UNSIGNED( 15 downto 0 );
      variable B : UNSIGNED( 15 downto 0 );
      variable Z : UNSIGNED( 0 downto 0 );
   begin
      A := ( dout_SegLenCnt_15_port, dout_SegLenCnt_14_port, 
            dout_SegLenCnt_13_port, dout_SegLenCnt_12_port, 
            dout_SegLenCnt_11_port, dout_SegLenCnt_10_port, 
            dout_SegLenCnt_9_port, dout_SegLenCnt_8_port, dout_SegLenCnt_7_port
            , dout_SegLenCnt_6_port, dout_SegLenCnt_5_port, 
            dout_SegLenCnt_4_port, dout_SegLenCnt_3_port, dout_SegLenCnt_2_port
            , dout_SegLenCnt_1_port, dout_SegLenCnt_0_port );
      B := ( X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port, X_Logic1_port, X_Logic0_port, X_Logic0_port );
      if ( A <= B ) then
         Z := ( others => '1' );
      else
         Z := ( others => '0' );
      end if;
      ( 0 => N40 ) <= Z;
   end process;
   
   eot_reg : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N170, next_state => cmd_25, 
               clocked_on => clk_port, Q => eot, QN => n_1150);
   decrypt_reg : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N182, next_state => cmd_28, 
               clocked_on => clk_port, Q => decrypt, QN => n_1151);
   bdoSIPO : DATA_SIPO_2 port map( clk => clk_port, rst => rst, end_of_input =>
                           end_of_block, data_p(31) => bdo_p_31_port, 
                           data_p(30) => bdo_p_30_port, data_p(29) => 
                           bdo_p_29_port, data_p(28) => bdo_p_28_port, 
                           data_p(27) => bdo_p_27_port, data_p(26) => 
                           bdo_p_26_port, data_p(25) => bdo_p_25_port, 
                           data_p(24) => bdo_p_24_port, data_p(23) => 
                           bdo_p_23_port, data_p(22) => bdo_p_22_port, 
                           data_p(21) => bdo_p_21_port, data_p(20) => 
                           bdo_p_20_port, data_p(19) => bdo_p_19_port, 
                           data_p(18) => bdo_p_18_port, data_p(17) => 
                           bdo_p_17_port, data_p(16) => bdo_p_16_port, 
                           data_p(15) => bdo_p_15_port, data_p(14) => 
                           bdo_p_14_port, data_p(13) => bdo_p_13_port, 
                           data_p(12) => bdo_p_12_port, data_p(11) => 
                           bdo_p_11_port, data_p(10) => bdo_p_10_port, 
                           data_p(9) => bdo_p_9_port, data_p(8) => bdo_p_8_port
                           , data_p(7) => bdo_p_7_port, data_p(6) => 
                           bdo_p_6_port, data_p(5) => bdo_p_5_port, data_p(4) 
                           => bdo_p_4_port, data_p(3) => bdo_p_3_port, 
                           data_p(2) => bdo_p_2_port, data_p(1) => bdo_p_1_port
                           , data_p(0) => bdo_p_0_port, data_valid_p => 
                           bdo_valid_p, data_ready_p => bdo_ready_p, data_s(31)
                           => bdo_cleared_31_port, data_s(30) => 
                           bdo_cleared_30_port, data_s(29) => 
                           bdo_cleared_29_port, data_s(28) => 
                           bdo_cleared_28_port, data_s(27) => 
                           bdo_cleared_27_port, data_s(26) => 
                           bdo_cleared_26_port, data_s(25) => 
                           bdo_cleared_25_port, data_s(24) => 
                           bdo_cleared_24_port, data_s(23) => 
                           bdo_cleared_23_port, data_s(22) => 
                           bdo_cleared_22_port, data_s(21) => 
                           bdo_cleared_21_port, data_s(20) => 
                           bdo_cleared_20_port, data_s(19) => 
                           bdo_cleared_19_port, data_s(18) => 
                           bdo_cleared_18_port, data_s(17) => 
                           bdo_cleared_17_port, data_s(16) => 
                           bdo_cleared_16_port, data_s(15) => 
                           bdo_cleared_15_port, data_s(14) => 
                           bdo_cleared_14_port, data_s(13) => 
                           bdo_cleared_13_port, data_s(12) => 
                           bdo_cleared_12_port, data_s(11) => 
                           bdo_cleared_11_port, data_s(10) => 
                           bdo_cleared_10_port, data_s(9) => bdo_cleared_9_port
                           , data_s(8) => bdo_cleared_8_port, data_s(7) => 
                           bdo_cleared_7_port, data_s(6) => bdo_cleared_6_port,
                           data_s(5) => bdo_cleared_5_port, data_s(4) => 
                           bdo_cleared_4_port, data_s(3) => bdo_cleared_3_port,
                           data_s(2) => bdo_cleared_2_port, data_s(1) => 
                           bdo_cleared_1_port, data_s(0) => bdo_cleared_0_port,
                           data_valid_s => bdo_valid, data_ready_s => bdo_ready
                           );
   pr_state_reg_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N184, next_state => N45, 
               clocked_on => clk_port, Q => pr_state_3_port, QN => n_1152);
   pr_state_reg_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N184, next_state => N44, 
               clocked_on => clk_port, Q => pr_state_2_port, QN => n_1153);
   pr_state_reg_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N184, next_state => N43, 
               clocked_on => clk_port, Q => pr_state_1_port, QN => n_1154);
   pr_state_reg_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N184, next_state => N42, 
               clocked_on => clk_port, Q => pr_state_0_port, QN => n_1155);
   C150 : GTECH_AND2 port map( A => N46, B => N47, Z => N50);
   C151 : GTECH_AND2 port map( A => N48, B => N49, Z => N51);
   C152 : GTECH_AND2 port map( A => N50, B => N51, Z => N52);
   C154 : GTECH_OR2 port map( A => pr_state_3_port, B => pr_state_2_port, Z => 
                           N53);
   C155 : GTECH_OR2 port map( A => pr_state_1_port, B => N49, Z => N54);
   C156 : GTECH_OR2 port map( A => N53, B => N54, Z => N55);
   C159 : GTECH_OR2 port map( A => pr_state_3_port, B => pr_state_2_port, Z => 
                           N57);
   C160 : GTECH_OR2 port map( A => N48, B => pr_state_0_port, Z => N58);
   C161 : GTECH_OR2 port map( A => N57, B => N58, Z => N59);
   C165 : GTECH_OR2 port map( A => pr_state_3_port, B => pr_state_2_port, Z => 
                           N61);
   C166 : GTECH_OR2 port map( A => N48, B => N49, Z => N62);
   C167 : GTECH_OR2 port map( A => N61, B => N62, Z => N63);
   C170 : GTECH_OR2 port map( A => pr_state_3_port, B => N47, Z => N65);
   C171 : GTECH_OR2 port map( A => pr_state_1_port, B => pr_state_0_port, Z => 
                           N66);
   C172 : GTECH_OR2 port map( A => N65, B => N66, Z => N67);
   C176 : GTECH_OR2 port map( A => pr_state_3_port, B => N47, Z => N69);
   C177 : GTECH_OR2 port map( A => pr_state_1_port, B => N49, Z => N70);
   C178 : GTECH_OR2 port map( A => N69, B => N70, Z => N71);
   C182 : GTECH_OR2 port map( A => pr_state_3_port, B => N47, Z => N73);
   C183 : GTECH_OR2 port map( A => N48, B => pr_state_0_port, Z => N74);
   C184 : GTECH_OR2 port map( A => N73, B => N74, Z => N75);
   C189 : GTECH_OR2 port map( A => pr_state_3_port, B => N47, Z => N77);
   C190 : GTECH_OR2 port map( A => N48, B => N49, Z => N78);
   C191 : GTECH_OR2 port map( A => N77, B => N78, Z => N79);
   C194 : GTECH_OR2 port map( A => N46, B => pr_state_2_port, Z => N81);
   C195 : GTECH_OR2 port map( A => pr_state_1_port, B => pr_state_0_port, Z => 
                           N82);
   C196 : GTECH_OR2 port map( A => N81, B => N82, Z => N83);
   C200 : GTECH_OR2 port map( A => N46, B => pr_state_2_port, Z => N85);
   C201 : GTECH_OR2 port map( A => pr_state_1_port, B => N49, Z => N86);
   C202 : GTECH_OR2 port map( A => N85, B => N86, Z => N87);
   C204 : GTECH_AND2 port map( A => pr_state_3_port, B => pr_state_1_port, Z =>
                           N89);
   C205 : GTECH_AND2 port map( A => pr_state_3_port, B => pr_state_2_port, Z =>
                           N90);
   C384 : GTECH_AND2 port map( A => N46, B => N47, Z => N116);
   C385 : GTECH_AND2 port map( A => N48, B => N49, Z => N117);
   C386 : GTECH_AND2 port map( A => N116, B => N117, Z => N118);
   C388 : GTECH_OR2 port map( A => pr_state_3_port, B => pr_state_2_port, Z => 
                           N119);
   C389 : GTECH_OR2 port map( A => pr_state_1_port, B => N49, Z => N120);
   C390 : GTECH_OR2 port map( A => N119, B => N120, Z => N121);
   C393 : GTECH_OR2 port map( A => pr_state_3_port, B => pr_state_2_port, Z => 
                           N123);
   C394 : GTECH_OR2 port map( A => N48, B => pr_state_0_port, Z => N124);
   C395 : GTECH_OR2 port map( A => N123, B => N124, Z => N125);
   C399 : GTECH_OR2 port map( A => pr_state_3_port, B => pr_state_2_port, Z => 
                           N127);
   C400 : GTECH_OR2 port map( A => N48, B => N49, Z => N128);
   C401 : GTECH_OR2 port map( A => N127, B => N128, Z => N129);
   C404 : GTECH_OR2 port map( A => pr_state_3_port, B => N47, Z => N131);
   C405 : GTECH_OR2 port map( A => pr_state_1_port, B => pr_state_0_port, Z => 
                           N132);
   C406 : GTECH_OR2 port map( A => N131, B => N132, Z => N133);
   C410 : GTECH_OR2 port map( A => pr_state_3_port, B => N47, Z => N135);
   C411 : GTECH_OR2 port map( A => pr_state_1_port, B => N49, Z => N136);
   C412 : GTECH_OR2 port map( A => N135, B => N136, Z => N137);
   C416 : GTECH_OR2 port map( A => pr_state_3_port, B => N47, Z => N139);
   C417 : GTECH_OR2 port map( A => N48, B => pr_state_0_port, Z => N140);
   C418 : GTECH_OR2 port map( A => N139, B => N140, Z => N141);
   C423 : GTECH_OR2 port map( A => pr_state_3_port, B => N47, Z => N143);
   C424 : GTECH_OR2 port map( A => N48, B => N49, Z => N144);
   C425 : GTECH_OR2 port map( A => N143, B => N144, Z => N145);
   C428 : GTECH_OR2 port map( A => N46, B => pr_state_2_port, Z => N147);
   C429 : GTECH_OR2 port map( A => pr_state_1_port, B => pr_state_0_port, Z => 
                           N148);
   C430 : GTECH_OR2 port map( A => N147, B => N148, Z => N149);
   C434 : GTECH_OR2 port map( A => N46, B => pr_state_2_port, Z => N151);
   C435 : GTECH_OR2 port map( A => pr_state_1_port, B => N49, Z => N152);
   C436 : GTECH_OR2 port map( A => N151, B => N152, Z => N153);
   C438 : GTECH_AND2 port map( A => pr_state_3_port, B => pr_state_1_port, Z =>
                           N155);
   C439 : GTECH_AND2 port map( A => pr_state_3_port, B => pr_state_2_port, Z =>
                           N156);
   I_0 : GTECH_NOT port map( A => cmd_31, Z => N185);
   C553 : GTECH_OR2 port map( A => cmd_30, B => N185, Z => N186);
   C554 : GTECH_OR2 port map( A => cmd_29, B => N186, Z => N187);
   C555 : GTECH_OR2 port map( A => cmd_28, B => N187, Z => N188);
   C557 : GTECH_OR2 port map( A => cmd_14_port, B => cmd_15_port, Z => N189);
   C558 : GTECH_OR2 port map( A => cmd_13_port, B => N189, Z => N190);
   C559 : GTECH_OR2 port map( A => cmd_12_port, B => N190, Z => N191);
   C560 : GTECH_OR2 port map( A => cmd_11_port, B => N191, Z => N192);
   C561 : GTECH_OR2 port map( A => cmd_10_port, B => N192, Z => N193);
   C562 : GTECH_OR2 port map( A => cmd_9_port, B => N193, Z => N194);
   C563 : GTECH_OR2 port map( A => cmd_8_port, B => N194, Z => N195);
   C564 : GTECH_OR2 port map( A => cmd_7_port, B => N195, Z => N196);
   C565 : GTECH_OR2 port map( A => cmd_6_port, B => N196, Z => N197);
   C566 : GTECH_OR2 port map( A => cmd_5_port, B => N197, Z => N198);
   C567 : GTECH_OR2 port map( A => cmd_4_port, B => N198, Z => N199);
   C568 : GTECH_OR2 port map( A => cmd_3_port, B => N199, Z => N200);
   C569 : GTECH_OR2 port map( A => cmd_2_port, B => N200, Z => N201);
   C570 : GTECH_OR2 port map( A => cmd_1_port, B => N201, Z => N202);
   C571 : GTECH_OR2 port map( A => cmd_0_port, B => N202, Z => N203);
   I_1 : GTECH_NOT port map( A => N203, Z => N204);
   C609_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 32 )
      port map(
         -- Connections to port 'DATA1'
         DATA(31) => do_data_internal_31_port, DATA(30) => 
               do_data_internal_30_port, DATA(29) => do_data_internal_29_port, 
               DATA(28) => do_data_internal_28_port, DATA(27) => 
               do_data_internal_27_port, DATA(26) => do_data_internal_26_port, 
               DATA(25) => do_data_internal_25_port, DATA(24) => 
               do_data_internal_24_port, DATA(23) => do_data_internal_23_port, 
               DATA(22) => do_data_internal_22_port, DATA(21) => 
               do_data_internal_21_port, DATA(20) => do_data_internal_20_port, 
               DATA(19) => do_data_internal_19_port, DATA(18) => 
               do_data_internal_18_port, DATA(17) => do_data_internal_17_port, 
               DATA(16) => do_data_internal_16_port, DATA(15) => 
               do_data_internal_15_port, DATA(14) => do_data_internal_14_port, 
               DATA(13) => do_data_internal_13_port, DATA(12) => 
               do_data_internal_12_port, DATA(11) => do_data_internal_11_port, 
               DATA(10) => do_data_internal_10_port, DATA(9) => 
               do_data_internal_9_port, DATA(8) => do_data_internal_8_port, 
               DATA(7) => do_data_internal_7_port, DATA(6) => 
               do_data_internal_6_port, DATA(5) => do_data_internal_5_port, 
               DATA(4) => do_data_internal_4_port, DATA(3) => 
               do_data_internal_3_port, DATA(2) => do_data_internal_2_port, 
               DATA(1) => do_data_internal_1_port, DATA(0) => 
               do_data_internal_0_port, 
         -- Connections to port 'DATA2'
         DATA(63) => X_Logic0_port, DATA(62) => X_Logic0_port, DATA(61) => 
               X_Logic0_port, DATA(60) => X_Logic0_port, DATA(59) => 
               X_Logic0_port, DATA(58) => X_Logic0_port, DATA(57) => 
               X_Logic0_port, DATA(56) => X_Logic0_port, DATA(55) => 
               X_Logic0_port, DATA(54) => X_Logic0_port, DATA(53) => 
               X_Logic0_port, DATA(52) => X_Logic0_port, DATA(51) => 
               X_Logic0_port, DATA(50) => X_Logic0_port, DATA(49) => 
               X_Logic0_port, DATA(48) => X_Logic0_port, DATA(47) => 
               X_Logic0_port, DATA(46) => X_Logic0_port, DATA(45) => 
               X_Logic0_port, DATA(44) => X_Logic0_port, DATA(43) => 
               X_Logic0_port, DATA(42) => X_Logic0_port, DATA(41) => 
               X_Logic0_port, DATA(40) => X_Logic0_port, DATA(39) => 
               X_Logic0_port, DATA(38) => X_Logic0_port, DATA(37) => 
               X_Logic0_port, DATA(36) => X_Logic0_port, DATA(35) => 
               X_Logic0_port, DATA(34) => X_Logic0_port, DATA(33) => 
               X_Logic0_port, DATA(32) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N0, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N1, 
         -- Connections to port 'Z'
         Z(31) => do_data_31_port, Z(30) => do_data_30_port, Z(29) => 
               do_data_29_port, Z(28) => do_data_28_port, Z(27) => 
               do_data_27_port, Z(26) => do_data_26_port, Z(25) => 
               do_data_25_port, Z(24) => do_data_24_port, Z(23) => 
               do_data_23_port, Z(22) => do_data_22_port, Z(21) => 
               do_data_21_port, Z(20) => do_data_20_port, Z(19) => 
               do_data_19_port, Z(18) => do_data_18_port, Z(17) => 
               do_data_17_port, Z(16) => do_data_16_port, Z(15) => 
               do_data_15_port, Z(14) => do_data_14_port, Z(13) => 
               do_data_13_port, Z(12) => do_data_12_port, Z(11) => 
               do_data_11_port, Z(10) => do_data_10_port, Z(9) => 
               do_data_9_port, Z(8) => do_data_8_port, Z(7) => do_data_7_port, 
               Z(6) => do_data_6_port, Z(5) => do_data_5_port, Z(4) => 
               do_data_4_port, Z(3) => do_data_3_port, Z(2) => do_data_2_port, 
               Z(1) => do_data_1_port, Z(0) => do_data_0_port );
   B_0 : GTECH_BUF port map( A => do_valid_port, Z => N0);
   B_1 : GTECH_BUF port map( A => N39, Z => N1);
   C610_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 4 )
      port map(
         -- Connections to port 'DATA1'
         DATA(3) => X_Logic0_port, DATA(2) => X_Logic0_port, DATA(1) => 
               X_Logic0_port, DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(7) => nx_state_3_port, DATA(6) => nx_state_2_port, DATA(5) => 
               nx_state_1_port, DATA(4) => nx_state_0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N2, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N3, 
         -- Connections to port 'Z'
         Z(3) => N45, Z(2) => N44, Z(1) => N43, Z(0) => N42 );
   B_2 : GTECH_BUF port map( A => rst, Z => N2);
   B_3 : GTECH_BUF port map( A => N41, Z => N3);
   C612_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => N188, 
         -- Connections to port 'DATA2'
         DATA(1) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N4, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N5, 
         -- Connections to port 'Z'
         Z(0) => N93 );
   B_4 : GTECH_BUF port map( A => cmd_valid_port, Z => N4);
   B_5 : GTECH_BUF port map( A => N92, Z => N5);
   I_2 : GTECH_NOT port map( A => N94, Z => N95);
   C614_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => decrypt, 
         -- Connections to port 'DATA2'
         DATA(1) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N6, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N7, 
         -- Connections to port 'Z'
         Z(0) => N98 );
   B_6 : GTECH_BUF port map( A => N204, Z => N6);
   B_7 : GTECH_BUF port map( A => N203, Z => N7);
   C615_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 2 )
      port map(
         -- Connections to port 'DATA1'
         DATA(1) => N98, DATA(0) => N204, 
         -- Connections to port 'DATA2'
         DATA(3) => X_Logic1_port, DATA(2) => X_Logic1_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N8, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N97, 
         -- Connections to port 'Z'
         Z(1) => N100, Z(0) => N99 );
   B_8 : GTECH_BUF port map( A => N96, Z => N8);
   C616_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => decrypt, 
         -- Connections to port 'DATA2'
         DATA(1) => X_Logic1_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N9, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N10, 
         -- Connections to port 'Z'
         Z(0) => N105 );
   B_9 : GTECH_BUF port map( A => eot, Z => N9);
   B_10 : GTECH_BUF port map( A => N104, Z => N10);
   C617_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 2 )
      port map(
         -- Connections to port 'DATA1'
         DATA(1) => eot, DATA(0) => N105, 
         -- Connections to port 'DATA2'
         DATA(3) => X_Logic1_port, DATA(2) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N11, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N12, 
         -- Connections to port 'Z'
         Z(1) => N107, Z(0) => N106 );
   B_11 : GTECH_BUF port map( A => last_flit_of_segment, Z => N11);
   B_12 : GTECH_BUF port map( A => N103, Z => N12);
   C618_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 3 )
      port map(
         -- Connections to port 'DATA1'
         DATA(2) => N107, DATA(1) => N106, DATA(0) => last_flit_of_segment, 
         -- Connections to port 'DATA2'
         DATA(5) => X_Logic1_port, DATA(4) => X_Logic0_port, DATA(3) => 
               X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N13, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N102, 
         -- Connections to port 'Z'
         Z(2) => N110, Z(1) => N109, Z(0) => N108 );
   B_13 : GTECH_BUF port map( A => N101, Z => N13);
   I_3 : GTECH_NOT port map( A => N111, Z => N112);
   C620_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => msg_auth_port, 
         -- Connections to port 'DATA2'
         DATA(1) => X_Logic1_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N14, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N15, 
         -- Connections to port 'Z'
         Z(0) => N114 );
   B_14 : GTECH_BUF port map( A => msg_auth_valid_port, Z => N14);
   B_15 : GTECH_BUF port map( A => N113, Z => N15);
   C621_cell : SELECT_OP
      generic map ( num_inputs => 10, input_width => 4 )
      port map(
         -- Connections to port 'DATA1'
         DATA(3) => X_Logic0_port, DATA(2) => X_Logic0_port, DATA(1) => N93, 
               DATA(0) => cmd_valid_port, 
         -- Connections to port 'DATA2'
         DATA(7) => X_Logic0_port, DATA(6) => X_Logic0_port, DATA(5) => 
               do_ready_port, DATA(4) => N115, 
         -- Connections to port 'DATA3'
         DATA(11) => N94, DATA(10) => X_Logic0_port, DATA(9) => N95, DATA(8) =>
               N94, 
         -- Connections to port 'DATA4'
         DATA(15) => X_Logic0_port, DATA(14) => N96, DATA(13) => N100, DATA(12)
               => N99, 
         -- Connections to port 'DATA5'
         DATA(19) => X_Logic0_port, DATA(18) => N110, DATA(17) => N109, 
               DATA(16) => N108, 
         -- Connections to port 'DATA6'
         DATA(23) => X_Logic0_port, DATA(22) => X_Logic1_port, DATA(21) => 
               do_ready_port, DATA(20) => N115, 
         -- Connections to port 'DATA7'
         DATA(27) => N111, DATA(26) => N112, DATA(25) => N112, DATA(24) => N111
               , 
         -- Connections to port 'DATA8'
         DATA(31) => msg_auth_valid_port, DATA(30) => N113, DATA(29) => N113, 
               DATA(28) => N114, 
         -- Connections to port 'DATA9'
         DATA(35) => N115, DATA(34) => X_Logic0_port, DATA(33) => X_Logic0_port
               , DATA(32) => X_Logic0_port, 
         -- Connections to port 'DATA10'
         DATA(39) => N115, DATA(38) => X_Logic0_port, DATA(37) => X_Logic0_port
               , DATA(36) => N115, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N16, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N17, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N18, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N19, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N20, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N21, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N22, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N23, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N24, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N25, 
         -- Connections to port 'Z'
         Z(3) => nx_state_3_port, Z(2) => nx_state_2_port, Z(1) => 
               nx_state_1_port, Z(0) => nx_state_0_port );
   B_16 : GTECH_BUF port map( A => N52, Z => N16);
   B_17 : GTECH_BUF port map( A => N56, Z => N17);
   B_18 : GTECH_BUF port map( A => N60, Z => N18);
   B_19 : GTECH_BUF port map( A => N64, Z => N19);
   B_20 : GTECH_BUF port map( A => N68, Z => N20);
   B_21 : GTECH_BUF port map( A => N72, Z => N21);
   B_22 : GTECH_BUF port map( A => N76, Z => N22);
   B_23 : GTECH_BUF port map( A => N80, Z => N23);
   B_24 : GTECH_BUF port map( A => N84, Z => N24);
   B_25 : GTECH_BUF port map( A => N88, Z => N25);
   C622_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => cmd_25, 
         -- Connections to port 'DATA2'
         DATA(1) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N26, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N27, 
         -- Connections to port 'Z'
         Z(0) => N160 );
   B_26 : GTECH_BUF port map( A => decrypt, Z => N26);
   B_27 : GTECH_BUF port map( A => N159, Z => N27);
   C623_cell : SELECT_OP
      generic map ( num_inputs => 11, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic1_port, 
         -- Connections to port 'DATA2'
         DATA(1) => X_Logic0_port, 
         -- Connections to port 'DATA3'
         DATA(2) => X_Logic0_port, 
         -- Connections to port 'DATA4'
         DATA(3) => do_ready_port, 
         -- Connections to port 'DATA5'
         DATA(4) => X_Logic0_port, 
         -- Connections to port 'DATA6'
         DATA(5) => X_Logic0_port, 
         -- Connections to port 'DATA7'
         DATA(6) => X_Logic0_port, 
         -- Connections to port 'DATA8'
         DATA(7) => X_Logic0_port, 
         -- Connections to port 'DATA9'
         DATA(8) => X_Logic0_port, 
         -- Connections to port 'DATA10'
         DATA(9) => X_Logic0_port, 
         -- Connections to port 'DATA11'
         DATA(10) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N28, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N29, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N30, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N31, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N32, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N33, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N34, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N35, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N36, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N37, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N38, 
         -- Connections to port 'Z'
         Z(0) => cmd_ready_port );
   B_28 : GTECH_BUF port map( A => N118, Z => N28);
   B_29 : GTECH_BUF port map( A => N122, Z => N29);
   B_30 : GTECH_BUF port map( A => N126, Z => N30);
   B_31 : GTECH_BUF port map( A => N130, Z => N31);
   B_32 : GTECH_BUF port map( A => N134, Z => N32);
   B_33 : GTECH_BUF port map( A => N138, Z => N33);
   B_34 : GTECH_BUF port map( A => N142, Z => N34);
   B_35 : GTECH_BUF port map( A => N146, Z => N35);
   B_36 : GTECH_BUF port map( A => N150, Z => N36);
   B_37 : GTECH_BUF port map( A => N154, Z => N37);
   B_38 : GTECH_BUF port map( A => N157, Z => N38);
   C624_cell : SELECT_OP
      generic map ( num_inputs => 11, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => X_Logic1_port, 
         -- Connections to port 'DATA3'
         DATA(2) => bdo_valid_p, 
         -- Connections to port 'DATA4'
         DATA(3) => cmd_valid_port, 
         -- Connections to port 'DATA5'
         DATA(4) => bdo_valid_p, 
         -- Connections to port 'DATA6'
         DATA(5) => X_Logic1_port, 
         -- Connections to port 'DATA7'
         DATA(6) => bdo_valid_p, 
         -- Connections to port 'DATA8'
         DATA(7) => X_Logic0_port, 
         -- Connections to port 'DATA9'
         DATA(8) => X_Logic1_port, 
         -- Connections to port 'DATA10'
         DATA(9) => X_Logic1_port, 
         -- Connections to port 'DATA11'
         DATA(10) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N28, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N29, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N30, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N31, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N32, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N33, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N34, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N35, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N36, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N37, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N38, 
         -- Connections to port 'Z'
         Z(0) => do_valid_port );
   C625_cell : SELECT_OP
      generic map ( num_inputs => 8, input_width => 32 )
      port map(
         -- Connections to port 'DATA1'
         DATA(31) => X_Logic1_port, DATA(30) => X_Logic0_port, DATA(29) => 
               X_Logic0_port, DATA(28) => X_Logic1_port, DATA(27) => 
               X_Logic0_port, DATA(26) => X_Logic0_port, DATA(25) => 
               X_Logic1_port, DATA(24) => X_Logic1_port, DATA(23) => 
               X_Logic0_port, DATA(22) => X_Logic0_port, DATA(21) => 
               X_Logic0_port, DATA(20) => X_Logic0_port, DATA(19) => 
               X_Logic0_port, DATA(18) => X_Logic0_port, DATA(17) => 
               X_Logic0_port, DATA(16) => X_Logic0_port, DATA(15) => 
               X_Logic0_port, DATA(14) => X_Logic0_port, DATA(13) => 
               X_Logic0_port, DATA(12) => X_Logic0_port, DATA(11) => 
               X_Logic0_port, DATA(10) => X_Logic0_port, DATA(9) => 
               X_Logic0_port, DATA(8) => X_Logic0_port, DATA(7) => 
               X_Logic0_port, DATA(6) => X_Logic0_port, DATA(5) => 
               X_Logic1_port, DATA(4) => X_Logic0_port, DATA(3) => 
               X_Logic0_port, DATA(2) => X_Logic0_port, DATA(1) => 
               X_Logic0_port, DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(63) => bdo_p_31_port, DATA(62) => bdo_p_30_port, DATA(61) => 
               bdo_p_29_port, DATA(60) => bdo_p_28_port, DATA(59) => 
               bdo_p_27_port, DATA(58) => bdo_p_26_port, DATA(57) => 
               bdo_p_25_port, DATA(56) => bdo_p_24_port, DATA(55) => 
               bdo_p_23_port, DATA(54) => bdo_p_22_port, DATA(53) => 
               bdo_p_21_port, DATA(52) => bdo_p_20_port, DATA(51) => 
               bdo_p_19_port, DATA(50) => bdo_p_18_port, DATA(49) => 
               bdo_p_17_port, DATA(48) => bdo_p_16_port, DATA(47) => 
               bdo_p_15_port, DATA(46) => bdo_p_14_port, DATA(45) => 
               bdo_p_13_port, DATA(44) => bdo_p_12_port, DATA(43) => 
               bdo_p_11_port, DATA(42) => bdo_p_10_port, DATA(41) => 
               bdo_p_9_port, DATA(40) => bdo_p_8_port, DATA(39) => bdo_p_7_port
               , DATA(38) => bdo_p_6_port, DATA(37) => bdo_p_5_port, DATA(36) 
               => bdo_p_4_port, DATA(35) => bdo_p_3_port, DATA(34) => 
               bdo_p_2_port, DATA(33) => bdo_p_1_port, DATA(32) => bdo_p_0_port
               , 
         -- Connections to port 'DATA3'
         DATA(95) => X_Logic0_port, DATA(94) => X_Logic1_port, DATA(93) => 
               X_Logic0_port, DATA(92) => N159, DATA(91) => X_Logic0_port, 
               DATA(90) => X_Logic0_port, DATA(89) => cmd_25, DATA(88) => N160,
               DATA(87) => X_Logic0_port, DATA(86) => X_Logic0_port, DATA(85) 
               => X_Logic0_port, DATA(84) => X_Logic0_port, DATA(83) => 
               X_Logic0_port, DATA(82) => X_Logic0_port, DATA(81) => 
               X_Logic0_port, DATA(80) => X_Logic0_port, DATA(79) => 
               cmd_15_port, DATA(78) => cmd_14_port, DATA(77) => cmd_13_port, 
               DATA(76) => cmd_12_port, DATA(75) => cmd_11_port, DATA(74) => 
               cmd_10_port, DATA(73) => cmd_9_port, DATA(72) => cmd_8_port, 
               DATA(71) => cmd_7_port, DATA(70) => cmd_6_port, DATA(69) => 
               cmd_5_port, DATA(68) => cmd_4_port, DATA(67) => cmd_3_port, 
               DATA(66) => cmd_2_port, DATA(65) => cmd_1_port, DATA(64) => 
               cmd_0_port, 
         -- Connections to port 'DATA4'
         DATA(127) => bdo_p_31_port, DATA(126) => bdo_p_30_port, DATA(125) => 
               bdo_p_29_port, DATA(124) => bdo_p_28_port, DATA(123) => 
               bdo_p_27_port, DATA(122) => bdo_p_26_port, DATA(121) => 
               bdo_p_25_port, DATA(120) => bdo_p_24_port, DATA(119) => 
               bdo_p_23_port, DATA(118) => bdo_p_22_port, DATA(117) => 
               bdo_p_21_port, DATA(116) => bdo_p_20_port, DATA(115) => 
               bdo_p_19_port, DATA(114) => bdo_p_18_port, DATA(113) => 
               bdo_p_17_port, DATA(112) => bdo_p_16_port, DATA(111) => 
               bdo_p_15_port, DATA(110) => bdo_p_14_port, DATA(109) => 
               bdo_p_13_port, DATA(108) => bdo_p_12_port, DATA(107) => 
               bdo_p_11_port, DATA(106) => bdo_p_10_port, DATA(105) => 
               bdo_p_9_port, DATA(104) => bdo_p_8_port, DATA(103) => 
               bdo_p_7_port, DATA(102) => bdo_p_6_port, DATA(101) => 
               bdo_p_5_port, DATA(100) => bdo_p_4_port, DATA(99) => 
               bdo_p_3_port, DATA(98) => bdo_p_2_port, DATA(97) => bdo_p_1_port
               , DATA(96) => bdo_p_0_port, 
         -- Connections to port 'DATA5'
         DATA(159) => X_Logic1_port, DATA(158) => X_Logic0_port, DATA(157) => 
               X_Logic0_port, DATA(156) => X_Logic0_port, DATA(155) => 
               X_Logic0_port, DATA(154) => X_Logic0_port, DATA(153) => 
               X_Logic1_port, DATA(152) => X_Logic1_port, DATA(151) => 
               X_Logic0_port, DATA(150) => X_Logic0_port, DATA(149) => 
               X_Logic0_port, DATA(148) => X_Logic0_port, DATA(147) => 
               X_Logic0_port, DATA(146) => X_Logic0_port, DATA(145) => 
               X_Logic0_port, DATA(144) => X_Logic0_port, DATA(143) => 
               X_Logic0_port, DATA(142) => X_Logic0_port, DATA(141) => 
               X_Logic0_port, DATA(140) => X_Logic0_port, DATA(139) => 
               X_Logic0_port, DATA(138) => X_Logic0_port, DATA(137) => 
               X_Logic0_port, DATA(136) => X_Logic0_port, DATA(135) => 
               X_Logic0_port, DATA(134) => X_Logic0_port, DATA(133) => 
               X_Logic0_port, DATA(132) => X_Logic1_port, DATA(131) => 
               X_Logic0_port, DATA(130) => X_Logic0_port, DATA(129) => 
               X_Logic0_port, DATA(128) => X_Logic0_port, 
         -- Connections to port 'DATA6'
         DATA(191) => bdo_p_31_port, DATA(190) => bdo_p_30_port, DATA(189) => 
               bdo_p_29_port, DATA(188) => bdo_p_28_port, DATA(187) => 
               bdo_p_27_port, DATA(186) => bdo_p_26_port, DATA(185) => 
               bdo_p_25_port, DATA(184) => bdo_p_24_port, DATA(183) => 
               bdo_p_23_port, DATA(182) => bdo_p_22_port, DATA(181) => 
               bdo_p_21_port, DATA(180) => bdo_p_20_port, DATA(179) => 
               bdo_p_19_port, DATA(178) => bdo_p_18_port, DATA(177) => 
               bdo_p_17_port, DATA(176) => bdo_p_16_port, DATA(175) => 
               bdo_p_15_port, DATA(174) => bdo_p_14_port, DATA(173) => 
               bdo_p_13_port, DATA(172) => bdo_p_12_port, DATA(171) => 
               bdo_p_11_port, DATA(170) => bdo_p_10_port, DATA(169) => 
               bdo_p_9_port, DATA(168) => bdo_p_8_port, DATA(167) => 
               bdo_p_7_port, DATA(166) => bdo_p_6_port, DATA(165) => 
               bdo_p_5_port, DATA(164) => bdo_p_4_port, DATA(163) => 
               bdo_p_3_port, DATA(162) => bdo_p_2_port, DATA(161) => 
               bdo_p_1_port, DATA(160) => bdo_p_0_port, 
         -- Connections to port 'DATA7'
         DATA(223) => X_Logic1_port, DATA(222) => X_Logic1_port, DATA(221) => 
               X_Logic1_port, DATA(220) => X_Logic1_port, DATA(219) => 
               X_Logic0_port, DATA(218) => X_Logic0_port, DATA(217) => 
               X_Logic0_port, DATA(216) => X_Logic0_port, DATA(215) => 
               X_Logic0_port, DATA(214) => X_Logic0_port, DATA(213) => 
               X_Logic0_port, DATA(212) => X_Logic0_port, DATA(211) => 
               X_Logic0_port, DATA(210) => X_Logic0_port, DATA(209) => 
               X_Logic0_port, DATA(208) => X_Logic0_port, DATA(207) => 
               X_Logic0_port, DATA(206) => X_Logic0_port, DATA(205) => 
               X_Logic0_port, DATA(204) => X_Logic0_port, DATA(203) => 
               X_Logic0_port, DATA(202) => X_Logic0_port, DATA(201) => 
               X_Logic0_port, DATA(200) => X_Logic0_port, DATA(199) => 
               X_Logic0_port, DATA(198) => X_Logic0_port, DATA(197) => 
               X_Logic0_port, DATA(196) => X_Logic0_port, DATA(195) => 
               X_Logic0_port, DATA(194) => X_Logic0_port, DATA(193) => 
               X_Logic0_port, DATA(192) => X_Logic0_port, 
         -- Connections to port 'DATA8'
         DATA(255) => X_Logic1_port, DATA(254) => X_Logic1_port, DATA(253) => 
               X_Logic1_port, DATA(252) => X_Logic0_port, DATA(251) => 
               X_Logic0_port, DATA(250) => X_Logic0_port, DATA(249) => 
               X_Logic0_port, DATA(248) => X_Logic0_port, DATA(247) => 
               X_Logic0_port, DATA(246) => X_Logic0_port, DATA(245) => 
               X_Logic0_port, DATA(244) => X_Logic0_port, DATA(243) => 
               X_Logic0_port, DATA(242) => X_Logic0_port, DATA(241) => 
               X_Logic0_port, DATA(240) => X_Logic0_port, DATA(239) => 
               X_Logic0_port, DATA(238) => X_Logic0_port, DATA(237) => 
               X_Logic0_port, DATA(236) => X_Logic0_port, DATA(235) => 
               X_Logic0_port, DATA(234) => X_Logic0_port, DATA(233) => 
               X_Logic0_port, DATA(232) => X_Logic0_port, DATA(231) => 
               X_Logic0_port, DATA(230) => X_Logic0_port, DATA(229) => 
               X_Logic0_port, DATA(228) => X_Logic0_port, DATA(227) => 
               X_Logic0_port, DATA(226) => X_Logic0_port, DATA(225) => 
               X_Logic0_port, DATA(224) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N29, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N30, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N31, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N32, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N33, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N34, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N36, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N37, 
         -- Connections to port 'Z'
         Z(31) => do_data_internal_31_port, Z(30) => do_data_internal_30_port, 
               Z(29) => do_data_internal_29_port, Z(28) => 
               do_data_internal_28_port, Z(27) => do_data_internal_27_port, 
               Z(26) => do_data_internal_26_port, Z(25) => 
               do_data_internal_25_port, Z(24) => do_data_internal_24_port, 
               Z(23) => do_data_internal_23_port, Z(22) => 
               do_data_internal_22_port, Z(21) => do_data_internal_21_port, 
               Z(20) => do_data_internal_20_port, Z(19) => 
               do_data_internal_19_port, Z(18) => do_data_internal_18_port, 
               Z(17) => do_data_internal_17_port, Z(16) => 
               do_data_internal_16_port, Z(15) => do_data_internal_15_port, 
               Z(14) => do_data_internal_14_port, Z(13) => 
               do_data_internal_13_port, Z(12) => do_data_internal_12_port, 
               Z(11) => do_data_internal_11_port, Z(10) => 
               do_data_internal_10_port, Z(9) => do_data_internal_9_port, Z(8) 
               => do_data_internal_8_port, Z(7) => do_data_internal_7_port, 
               Z(6) => do_data_internal_6_port, Z(5) => do_data_internal_5_port
               , Z(4) => do_data_internal_4_port, Z(3) => 
               do_data_internal_3_port, Z(2) => do_data_internal_2_port, Z(1) 
               => do_data_internal_1_port, Z(0) => do_data_internal_0_port );
   C626_cell : SELECT_OP
      generic map ( num_inputs => 11, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => X_Logic0_port, 
         -- Connections to port 'DATA3'
         DATA(2) => do_ready_port, 
         -- Connections to port 'DATA4'
         DATA(3) => X_Logic0_port, 
         -- Connections to port 'DATA5'
         DATA(4) => do_ready_port, 
         -- Connections to port 'DATA6'
         DATA(5) => X_Logic0_port, 
         -- Connections to port 'DATA7'
         DATA(6) => do_ready_port, 
         -- Connections to port 'DATA8'
         DATA(7) => X_Logic0_port, 
         -- Connections to port 'DATA9'
         DATA(8) => X_Logic0_port, 
         -- Connections to port 'DATA10'
         DATA(9) => X_Logic0_port, 
         -- Connections to port 'DATA11'
         DATA(10) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N28, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N29, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N30, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N31, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N32, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N33, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N34, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N35, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N36, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N37, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N38, 
         -- Connections to port 'Z'
         Z(0) => bdo_ready_p );
   C627_cell : SELECT_OP
      generic map ( num_inputs => 11, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => X_Logic0_port, 
         -- Connections to port 'DATA3'
         DATA(2) => X_Logic0_port, 
         -- Connections to port 'DATA4'
         DATA(3) => N158, 
         -- Connections to port 'DATA5'
         DATA(4) => X_Logic0_port, 
         -- Connections to port 'DATA6'
         DATA(5) => X_Logic0_port, 
         -- Connections to port 'DATA7'
         DATA(6) => X_Logic0_port, 
         -- Connections to port 'DATA8'
         DATA(7) => X_Logic0_port, 
         -- Connections to port 'DATA9'
         DATA(8) => X_Logic0_port, 
         -- Connections to port 'DATA10'
         DATA(9) => X_Logic0_port, 
         -- Connections to port 'DATA11'
         DATA(10) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N28, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N29, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N30, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N31, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N32, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N33, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N34, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N35, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N36, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N37, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N38, 
         -- Connections to port 'Z'
         Z(0) => len_SegLenCnt );
   C628_cell : SELECT_OP
      generic map ( num_inputs => 11, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => X_Logic0_port, 
         -- Connections to port 'DATA3'
         DATA(2) => X_Logic0_port, 
         -- Connections to port 'DATA4'
         DATA(3) => X_Logic0_port, 
         -- Connections to port 'DATA5'
         DATA(4) => N101, 
         -- Connections to port 'DATA6'
         DATA(5) => X_Logic0_port, 
         -- Connections to port 'DATA7'
         DATA(6) => X_Logic0_port, 
         -- Connections to port 'DATA8'
         DATA(7) => X_Logic0_port, 
         -- Connections to port 'DATA9'
         DATA(8) => X_Logic0_port, 
         -- Connections to port 'DATA10'
         DATA(9) => X_Logic0_port, 
         -- Connections to port 'DATA11'
         DATA(10) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N28, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N29, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N30, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N31, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N32, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N33, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N34, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N35, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N36, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N37, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N38, 
         -- Connections to port 'Z'
         Z(0) => en_SegLenCnt );
   C629_cell : SELECT_OP
      generic map ( num_inputs => 11, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => X_Logic0_port, 
         -- Connections to port 'DATA3'
         DATA(2) => X_Logic0_port, 
         -- Connections to port 'DATA4'
         DATA(3) => X_Logic0_port, 
         -- Connections to port 'DATA5'
         DATA(4) => X_Logic0_port, 
         -- Connections to port 'DATA6'
         DATA(5) => X_Logic0_port, 
         -- Connections to port 'DATA7'
         DATA(6) => X_Logic0_port, 
         -- Connections to port 'DATA8'
         DATA(7) => X_Logic1_port, 
         -- Connections to port 'DATA9'
         DATA(8) => X_Logic0_port, 
         -- Connections to port 'DATA10'
         DATA(9) => X_Logic0_port, 
         -- Connections to port 'DATA11'
         DATA(10) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N28, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N29, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N30, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N31, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N32, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N33, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N34, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N35, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N36, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N37, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N38, 
         -- Connections to port 'Z'
         Z(0) => msg_auth_ready_port );
   C630_cell : SELECT_OP
      generic map ( num_inputs => 11, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => X_Logic0_port, 
         -- Connections to port 'DATA3'
         DATA(2) => X_Logic0_port, 
         -- Connections to port 'DATA4'
         DATA(3) => X_Logic0_port, 
         -- Connections to port 'DATA5'
         DATA(4) => X_Logic0_port, 
         -- Connections to port 'DATA6'
         DATA(5) => X_Logic0_port, 
         -- Connections to port 'DATA7'
         DATA(6) => X_Logic0_port, 
         -- Connections to port 'DATA8'
         DATA(7) => X_Logic0_port, 
         -- Connections to port 'DATA9'
         DATA(8) => X_Logic1_port, 
         -- Connections to port 'DATA10'
         DATA(9) => X_Logic1_port, 
         -- Connections to port 'DATA11'
         DATA(10) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N28, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N29, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N30, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N31, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N32, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N33, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N34, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N35, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N36, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N37, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N38, 
         -- Connections to port 'Z'
         Z(0) => do_last_port );
         X_Logic1_port <= '1';
         X_Logic0_port <= '0';
   C637 : GTECH_AND2 port map( A => bdo(31), B => bdo_valid_bytes(3), Z => 
                           bdo_cleared_31_port);
   C638 : GTECH_AND2 port map( A => bdo(30), B => bdo_valid_bytes(3), Z => 
                           bdo_cleared_30_port);
   C639 : GTECH_AND2 port map( A => bdo(29), B => bdo_valid_bytes(3), Z => 
                           bdo_cleared_29_port);
   C640 : GTECH_AND2 port map( A => bdo(28), B => bdo_valid_bytes(3), Z => 
                           bdo_cleared_28_port);
   C641 : GTECH_AND2 port map( A => bdo(27), B => bdo_valid_bytes(3), Z => 
                           bdo_cleared_27_port);
   C642 : GTECH_AND2 port map( A => bdo(26), B => bdo_valid_bytes(3), Z => 
                           bdo_cleared_26_port);
   C643 : GTECH_AND2 port map( A => bdo(25), B => bdo_valid_bytes(3), Z => 
                           bdo_cleared_25_port);
   C644 : GTECH_AND2 port map( A => bdo(24), B => bdo_valid_bytes(3), Z => 
                           bdo_cleared_24_port);
   C645 : GTECH_AND2 port map( A => bdo(23), B => bdo_valid_bytes(2), Z => 
                           bdo_cleared_23_port);
   C646 : GTECH_AND2 port map( A => bdo(22), B => bdo_valid_bytes(2), Z => 
                           bdo_cleared_22_port);
   C647 : GTECH_AND2 port map( A => bdo(21), B => bdo_valid_bytes(2), Z => 
                           bdo_cleared_21_port);
   C648 : GTECH_AND2 port map( A => bdo(20), B => bdo_valid_bytes(2), Z => 
                           bdo_cleared_20_port);
   C649 : GTECH_AND2 port map( A => bdo(19), B => bdo_valid_bytes(2), Z => 
                           bdo_cleared_19_port);
   C650 : GTECH_AND2 port map( A => bdo(18), B => bdo_valid_bytes(2), Z => 
                           bdo_cleared_18_port);
   C651 : GTECH_AND2 port map( A => bdo(17), B => bdo_valid_bytes(2), Z => 
                           bdo_cleared_17_port);
   C652 : GTECH_AND2 port map( A => bdo(16), B => bdo_valid_bytes(2), Z => 
                           bdo_cleared_16_port);
   C653 : GTECH_AND2 port map( A => bdo(15), B => bdo_valid_bytes(1), Z => 
                           bdo_cleared_15_port);
   C654 : GTECH_AND2 port map( A => bdo(14), B => bdo_valid_bytes(1), Z => 
                           bdo_cleared_14_port);
   C655 : GTECH_AND2 port map( A => bdo(13), B => bdo_valid_bytes(1), Z => 
                           bdo_cleared_13_port);
   C656 : GTECH_AND2 port map( A => bdo(12), B => bdo_valid_bytes(1), Z => 
                           bdo_cleared_12_port);
   C657 : GTECH_AND2 port map( A => bdo(11), B => bdo_valid_bytes(1), Z => 
                           bdo_cleared_11_port);
   C658 : GTECH_AND2 port map( A => bdo(10), B => bdo_valid_bytes(1), Z => 
                           bdo_cleared_10_port);
   C659 : GTECH_AND2 port map( A => bdo(9), B => bdo_valid_bytes(1), Z => 
                           bdo_cleared_9_port);
   C660 : GTECH_AND2 port map( A => bdo(8), B => bdo_valid_bytes(1), Z => 
                           bdo_cleared_8_port);
   C661 : GTECH_AND2 port map( A => bdo(7), B => bdo_valid_bytes(0), Z => 
                           bdo_cleared_7_port);
   C662 : GTECH_AND2 port map( A => bdo(6), B => bdo_valid_bytes(0), Z => 
                           bdo_cleared_6_port);
   C663 : GTECH_AND2 port map( A => bdo(5), B => bdo_valid_bytes(0), Z => 
                           bdo_cleared_5_port);
   C664 : GTECH_AND2 port map( A => bdo(4), B => bdo_valid_bytes(0), Z => 
                           bdo_cleared_4_port);
   C665 : GTECH_AND2 port map( A => bdo(3), B => bdo_valid_bytes(0), Z => 
                           bdo_cleared_3_port);
   C666 : GTECH_AND2 port map( A => bdo(2), B => bdo_valid_bytes(0), Z => 
                           bdo_cleared_2_port);
   C667 : GTECH_AND2 port map( A => bdo(1), B => bdo_valid_bytes(0), Z => 
                           bdo_cleared_1_port);
   C668 : GTECH_AND2 port map( A => bdo(0), B => bdo_valid_bytes(0), Z => 
                           bdo_cleared_0_port);
   I_4 : GTECH_NOT port map( A => do_valid_port, Z => N39);
   B_39 : GTECH_BUF port map( A => N40, Z => last_flit_of_segment);
   I_5 : GTECH_NOT port map( A => rst, Z => N41);
   I_6 : GTECH_NOT port map( A => pr_state_3_port, Z => N46);
   I_7 : GTECH_NOT port map( A => pr_state_2_port, Z => N47);
   I_8 : GTECH_NOT port map( A => pr_state_1_port, Z => N48);
   I_9 : GTECH_NOT port map( A => pr_state_0_port, Z => N49);
   I_10 : GTECH_NOT port map( A => N55, Z => N56);
   I_11 : GTECH_NOT port map( A => N59, Z => N60);
   I_12 : GTECH_NOT port map( A => N63, Z => N64);
   I_13 : GTECH_NOT port map( A => N67, Z => N68);
   I_14 : GTECH_NOT port map( A => N71, Z => N72);
   I_15 : GTECH_NOT port map( A => N75, Z => N76);
   I_16 : GTECH_NOT port map( A => N79, Z => N80);
   I_17 : GTECH_NOT port map( A => N83, Z => N84);
   I_18 : GTECH_NOT port map( A => N87, Z => N88);
   C704 : GTECH_OR2 port map( A => N89, B => N90, Z => N91);
   I_19 : GTECH_NOT port map( A => cmd_valid_port, Z => N92);
   C720 : GTECH_AND2 port map( A => N205, B => end_of_block, Z => N94);
   C721 : GTECH_AND2 port map( A => bdo_valid_p, B => do_ready_port, Z => N205)
                           ;
   C723 : GTECH_AND2 port map( A => cmd_valid_port, B => do_ready_port, Z => 
                           N96);
   I_20 : GTECH_NOT port map( A => N96, Z => N97);
   C729 : GTECH_AND2 port map( A => bdo_valid_p, B => do_ready_port, Z => N101)
                           ;
   I_21 : GTECH_NOT port map( A => N101, Z => N102);
   I_22 : GTECH_NOT port map( A => last_flit_of_segment, Z => N103);
   I_23 : GTECH_NOT port map( A => eot, Z => N104);
   C739 : GTECH_AND2 port map( A => N206, B => do_ready_port, Z => N111);
   C740 : GTECH_AND2 port map( A => bdo_valid_p, B => end_of_block, Z => N206);
   I_24 : GTECH_NOT port map( A => msg_auth_valid_port, Z => N113);
   I_25 : GTECH_NOT port map( A => do_ready_port, Z => N115);
   I_26 : GTECH_NOT port map( A => N121, Z => N122);
   I_27 : GTECH_NOT port map( A => N125, Z => N126);
   I_28 : GTECH_NOT port map( A => N129, Z => N130);
   I_29 : GTECH_NOT port map( A => N133, Z => N134);
   I_30 : GTECH_NOT port map( A => N137, Z => N138);
   I_31 : GTECH_NOT port map( A => N141, Z => N142);
   I_32 : GTECH_NOT port map( A => N145, Z => N146);
   I_33 : GTECH_NOT port map( A => N149, Z => N150);
   I_34 : GTECH_NOT port map( A => N153, Z => N154);
   C777 : GTECH_OR2 port map( A => N155, B => N156, Z => N157);
   C789 : GTECH_AND2 port map( A => do_ready_port, B => cmd_valid_port, Z => 
                           N158);
   I_35 : GTECH_NOT port map( A => decrypt, Z => N159);
   C793 : GTECH_OR2 port map( A => N118, B => N122, Z => N161);
   C794 : GTECH_OR2 port map( A => N161, B => N126, Z => N162);
   C795 : GTECH_OR2 port map( A => N162, B => N134, Z => N163);
   C796 : GTECH_OR2 port map( A => N163, B => N138, Z => N164);
   C797 : GTECH_OR2 port map( A => N164, B => N142, Z => N165);
   C798 : GTECH_OR2 port map( A => N165, B => N146, Z => N166);
   C799 : GTECH_OR2 port map( A => N166, B => N150, Z => N167);
   C800 : GTECH_OR2 port map( A => N167, B => N154, Z => N168);
   C801 : GTECH_OR2 port map( A => N168, B => N157, Z => N169);
   I_36 : GTECH_NOT port map( A => N169, Z => N170);
   C803 : GTECH_AND2 port map( A => N92, B => N118, Z => N171);
   C804 : GTECH_OR2 port map( A => N171, B => N122, Z => N172);
   C805 : GTECH_OR2 port map( A => N172, B => N126, Z => N173);
   C806 : GTECH_OR2 port map( A => N173, B => N130, Z => N174);
   C807 : GTECH_OR2 port map( A => N174, B => N134, Z => N175);
   C808 : GTECH_OR2 port map( A => N175, B => N138, Z => N176);
   C809 : GTECH_OR2 port map( A => N176, B => N142, Z => N177);
   C810 : GTECH_OR2 port map( A => N177, B => N146, Z => N178);
   C811 : GTECH_OR2 port map( A => N178, B => N150, Z => N179);
   C812 : GTECH_OR2 port map( A => N179, B => N154, Z => N180);
   C813 : GTECH_OR2 port map( A => N180, B => N157, Z => N181);
   I_37 : GTECH_NOT port map( A => N181, Z => N182);
   C815 : GTECH_AND2 port map( A => N91, B => N41, Z => N183);
   I_38 : GTECH_NOT port map( A => N183, Z => N184);

end SYN_PostProcessor;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_LWC_1.all;

entity CryptoCore_2 is

   port( clk, rst : in std_logic;  key : in std_logic_vector (31 downto 0);  
         key_valid : in std_logic;  key_ready : out std_logic;  bdi : in 
         std_logic_vector (31 downto 0);  bdi_valid : in std_logic;  bdi_ready 
         : out std_logic;  bdi_pad_loc, bdi_valid_bytes : in std_logic_vector 
         (3 downto 0);  bdi_size : in std_logic_vector (2 downto 0);  bdi_eot, 
         bdi_eoi : in std_logic;  bdi_type : in std_logic_vector (3 downto 0); 
         decrypt_in, key_update, hash_in : in std_logic;  bdo : out 
         std_logic_vector (31 downto 0);  bdo_valid : out std_logic;  bdo_ready
         : in std_logic;  bdo_type, bdo_valid_bytes : out std_logic_vector (3 
         downto 0);  end_of_block, msg_auth_valid : out std_logic;  
         msg_auth_ready : in std_logic;  msg_auth : out std_logic);

end CryptoCore_2;

architecture SYN_behavioral of CryptoCore_2 is

   component GTECH_NOT
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component GTECH_OR2
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component GTECH_AND2
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component GTECH_BUF
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
      generic ( ac_as_q, ac_as_qn, sc_ss_q : integer );
      port(
         clear, preset, enable, data_in, synch_clear, synch_preset, 
            synch_toggle, synch_enable, next_state, clocked_on : in std_logic;
         Q, QN : buffer std_logic
      );
   end component;
   
   component cyclist_ops_DATA_LEN32_1
      port( clk, key_en : in std_logic;  state_main_en : in std_logic_vector (2
            downto 0);  state_main_sel : in std_logic_vector (6 downto 0);  
            cyc_state_update_sel, xor_sel : in std_logic;  cycd_sel : in 
            std_logic_vector (1 downto 0);  extract_sel : in std_logic;  
            bdi_key : in std_logic_vector (31 downto 0);  cu_cd : in 
            std_logic_vector (7 downto 0);  dcount_in, rnd_counter : in 
            std_logic_vector (3 downto 0);  bdo_out : out std_logic_vector (31 
            downto 0));
   end component;
   
   component counter_num_bits4_1
      port( clk, reset, enable : in std_logic;  q : out std_logic_vector (3 
            downto 0));
   end component;
   
   signal N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15,
      N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30
      , N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, 
      N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59
      , N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N73, 
      N74, N75, X_Logic1_port, X_Logic0_port, clk_port, key_31_port, 
      key_30_port, key_29_port, key_28_port, key_27_port, key_26_port, 
      key_25_port, key_24_port, key_23_port, key_22_port, key_21_port, 
      key_20_port, key_19_port, key_18_port, key_17_port, key_16_port, 
      key_15_port, key_14_port, key_13_port, key_12_port, key_11_port, 
      key_10_port, key_9_port, key_8_port, key_7_port, key_6_port, key_5_port, 
      key_4_port, key_3_port, key_2_port, key_1_port, key_0_port, 
      key_valid_port, key_ready_port, bdi_31_port, bdi_30_port, bdi_29_port, 
      bdi_28_port, bdi_27_port, bdi_26_port, bdi_25_port, bdi_24_port, 
      bdi_23_port, bdi_22_port, bdi_21_port, bdi_20_port, bdi_19_port, 
      bdi_18_port, bdi_17_port, bdi_16_port, bdi_15_port, bdi_14_port, 
      bdi_13_port, bdi_12_port, bdi_11_port, bdi_10_port, bdi_9_port, 
      bdi_8_port, bdi_7_port, bdi_6_port, bdi_5_port, bdi_4_port, bdi_3_port, 
      bdi_2_port, bdi_1_port, bdi_0_port, bdi_valid_port, bdi_ready_port, 
      bdi_valid_bytes_3_port, bdi_valid_bytes_2_port, bdi_valid_bytes_1_port, 
      bdi_valid_bytes_0_port, bdi_size_2_port, bdi_size_1_port, bdi_size_0_port
      , bdi_eot_port, decrypt_in_port, key_update_port, hash_in_port, 
      bdo_31_port, bdo_30_port, bdo_29_port, bdo_28_port, bdo_27_port, 
      bdo_26_port, bdo_25_port, bdo_24_port, bdo_23_port, bdo_22_port, 
      bdo_21_port, bdo_20_port, bdo_19_port, bdo_18_port, bdo_17_port, 
      bdo_16_port, bdo_15_port, bdo_14_port, bdo_13_port, bdo_12_port, 
      bdo_11_port, bdo_10_port, bdo_9_port, bdo_8_port, bdo_7_port, bdo_6_port,
      bdo_5_port, bdo_4_port, bdo_3_port, bdo_2_port, bdo_1_port, bdo_0_port, 
      bdo_valid_port, bdo_ready_port, bdo_type_3_port, bdo_type_2_port, 
      bdo_type_0, bdo_valid_bytes_3_port, bdo_valid_bytes_2_port, 
      bdo_valid_bytes_1_port, bdo_valid_bytes_0_port, end_of_block_port, 
      msg_auth_valid_port, msg_auth_port, load_rnd, en_rnd, rnd_counter_3_port,
      rnd_counter_2_port, rnd_counter_1_port, rnd_counter_0_port, load_dcount, 
      en_dcount, dcount_3_port, dcount_2_port, dcount_1_port, dcount_0_port, 
      key_en, state_main_en_2_port, state_main_en_1_port, state_main_en_0_port,
      state_main_sel_6_port, state_main_sel_5_port, state_main_sel_4_port, 
      state_main_sel_2, state_main_sel_0, cyc_state_update_sel, xor_sel, 
      cycd_sel_1_port, cycd_sel_0_port, extract_sel, bdi_key_31_port, 
      bdi_key_30_port, bdi_key_29_port, bdi_key_28_port, bdi_key_27_port, 
      bdi_key_26_port, bdi_key_25_port, bdi_key_24_port, bdi_key_23_port, 
      bdi_key_22_port, bdi_key_21_port, bdi_key_20_port, bdi_key_19_port, 
      bdi_key_18_port, bdi_key_17_port, bdi_key_16_port, bdi_key_15_port, 
      bdi_key_14_port, bdi_key_13_port, bdi_key_12_port, bdi_key_11_port, 
      bdi_key_10_port, bdi_key_9_port, bdi_key_8_port, bdi_key_7_port, 
      bdi_key_6_port, bdi_key_5_port, bdi_key_4_port, bdi_key_3_port, 
      bdi_key_2_port, bdi_key_1_port, bdi_key_0_port, cu_cd_s_7_port, 
      cu_cd_s_6_port, cu_cd_s_1, cu_cd_s_0, cyc_s_2_port, cyc_s_1_port, 
      cyc_s_0_port, n_calling_state_2_port, n_calling_state_1_port, 
      n_calling_state_0_port, calling_state_2_port, calling_state_1_port, 
      calling_state_0_port, n_cyc_s_2_port, n_cyc_s_1_port, n_cyc_s_0_port, 
      mode_1_port, mode_0_port, n_decrypt_op_s, decrypt_op_s, n_tag_verified, 
      n_gtr_one_perm, gtr_one_perm, n_bdi_eot_prev, N76, N77, N78, N79, N80, 
      N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95
      , N96, N97, N98, N99, N100, N101, N102, N103, N104, N105, N106, N107, 
      N108, N109, N110, N111, N112, N113, N114, N115, N116, N117, N118, N119, 
      N120, N121, N122, N123, N124, N125, N126, N127, N128, N129, N130, N131, 
      N132, N133, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143, 
      N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154, N155, 
      N156, N157, N158, N159, N160, N161, N162, N163, N164, N165, N166, N167, 
      N168, N169, N170, N171, N172, N173, N174, N175, N176, N177, N178, N179, 
      N180, N181, N182, N183, N184, N185, N186, N187, N188, N189, N190, N191, 
      N192, N193, N194, N195, N196, N197, N198, N199, N200, N201, N202, N203, 
      N204, N205, N206, N207, N208, N209, N210, N211, N212, N213, N214, N215, 
      N216, N217, N218, N219, N220, N221, N222, N223, N224, N225, N226, N227, 
      N228, N229, N230, N231, N232, N233, N234, N235, N236, N237, N238, N239, 
      N240, N241, N242, N243, N244, N245, N246, N247, N248, N249, N250, N251, 
      N252, N253, N254, N255, N256, N257, N258, N259, N260, N261, N262, N263, 
      N264, N265, N266, N267, N268, N269, N270, N271, N272, N273, N274, N275, 
      N276, N277, N278, N279, N280, N281, N282, N283, N284, N285, N286, N287, 
      N288, N289, N290, N291, N292, N293, N294, N295, N296, N297, N298, N299, 
      N300, N301, N302, N303, N304, N305, N306, N307, N308, N309, N310, N311, 
      N312, N313, N314, N315, N316, N317, bdi_eot_prev, N318, N319, N320, N321,
      N322, N323, N324, N325, N326, N327, N328, N329, N330, N331, N332, N333, 
      N334, N335, N336, N337, N338, N339, N340, N341, N342, N343, N344, N345, 
      N346, N347, N348, N349, N350, N351, N352, N353, N354, N355, N356, N357, 
      N358, N359, N360, N361, N362, N363, N364, N365, N366, N367, N368, N369, 
      N370, N371, N372, N373, N374, N375, N376, N377, N378, N379, N380, N381, 
      N382, N383, N384, N385, N386, N387, N388, N389, N390, N391, N392, N393, 
      N394, N395, N396, N397, N398, N399, N400, N401, N402, N403, N404, N405, 
      N406, N407, N408, N409, N410, N411, N412, N413, N414, N415, N416, N417, 
      N418, N419, N420, N421, N422, N423, N424, N425, N426, N427, N428, N429, 
      N430, N431, N432, N433, N434, N435, N436, N437, N438, N439, N440, N441, 
      N442, N443, N444, N445, N446, N447, N448, N449, N450, N451, N452, N453, 
      N454, N455, N456, N457, N458, N459, N460, N461, N462, N463, N464, N465, 
      N466, N467, N468, N469, N470, N471, N472, N473, N474, N475, N476, N477, 
      N478, N479, N480, N481, N482, N483, N484, N485, N486, N487, N488, N489, 
      N490, N491, N492, N493, N494, N495, N496, N497, N498, N499, N500, N501, 
      N502, N503, N504, N505, N506, N507, N508, N509, N510, N511, N512, N513, 
      N514, N515, N516, N517, N518, N519, N520, N521, N522, N523, N524, N525, 
      N526, N527, N528, N529, N530, N531, N532, N533, N534, N535, N536, N537, 
      N538, N539, N540, N541, N542, N543, N544, N545, N546, N547, tag_verified,
      N548, N549, N550, N551, N552, N553, N554, N555, N556, N557, N558, N559, 
      N560, N561, N562, N563, N564, N565, N566, N567, N568, N569, N570, N571, 
      N572, N573, N574, N575, N576, N577, N578, N579, N580, N581, N582, N583, 
      N584, N585, N586, N587, N588, N589, N590, N591, N592, N593, N594, N595, 
      N596, N597, N598, N599, N600, N601, N602, N603, N604, N605, N606, N607, 
      N608, N609, N610, N611, N612, N613, N614, N615, N616, N617, N618, N619, 
      N620, N621, N622, N623, N624, N625, N626, N627, N628, N629, N630, N631, 
      N632, N633, N634, N635, N636, N637, N638, N639, N640, N641, N642, N643, 
      N644, N645, N646, N647, N648, N649, N650, N651, N652, N653, N654, N655, 
      N656, N657, N658, N659, N660, N661, N662, N663, N664, N665, N666, N667, 
      N668, N669, N670, N671, N672, N673, N674, N675, N676, N677, N678, N679, 
      N680, N681, N682, N683, N684, N685, N686, N687, N688, N689, N690, N691, 
      N692, N693, N694, N695, N696, N697, N698, N699, N700, N701, N702, N703, 
      N704, N705, N706, N707, N708, N709, N710, N711, N712, N713, N714, N715, 
      N716, N717, N718, N719, N720, N721, N722, N723, N724, N725, N726, N727, 
      N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, 
      N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, 
      N752, N753, N754, N755, N756, N757, N758, N759, N760, N761, N762, N763, 
      N764, N765, N766, N767, N768, N769, N770, N771, N772, N773, N774, N775, 
      N776, N777, N778, N779, N780, N781, N782, N783, N784, N785, N786, N787, 
      N788, N789, N790, N791, N792, N793, N794, N795, N796, N797, N798, N799, 
      N800, N801, N802, N803, N804, N805, N806, N807, N808, n_1156, n_1157, 
      n_1158, n_1159, n_1160, n_1161, n_1162, n_1163, n_1164, n_1165, n_1166, 
      n_1167, n_1168, n_1169, n_1170, n_1171, n_1172, n_1173, n_1174, n_1175, 
      n_1176, n_1177, n_1178 : std_logic;

begin
   clk_port <= clk;
   ( key_31_port, key_30_port, key_29_port, key_28_port, key_27_port, 
      key_26_port, key_25_port, key_24_port, key_23_port, key_22_port, 
      key_21_port, key_20_port, key_19_port, key_18_port, key_17_port, 
      key_16_port, key_15_port, key_14_port, key_13_port, key_12_port, 
      key_11_port, key_10_port, key_9_port, key_8_port, key_7_port, key_6_port,
      key_5_port, key_4_port, key_3_port, key_2_port, key_1_port, key_0_port ) 
      <= key;
   key_valid_port <= key_valid;
   key_ready <= key_ready_port;
   ( bdi_31_port, bdi_30_port, bdi_29_port, bdi_28_port, bdi_27_port, 
      bdi_26_port, bdi_25_port, bdi_24_port, bdi_23_port, bdi_22_port, 
      bdi_21_port, bdi_20_port, bdi_19_port, bdi_18_port, bdi_17_port, 
      bdi_16_port, bdi_15_port, bdi_14_port, bdi_13_port, bdi_12_port, 
      bdi_11_port, bdi_10_port, bdi_9_port, bdi_8_port, bdi_7_port, bdi_6_port,
      bdi_5_port, bdi_4_port, bdi_3_port, bdi_2_port, bdi_1_port, bdi_0_port ) 
      <= bdi;
   bdi_valid_port <= bdi_valid;
   bdi_ready <= bdi_ready_port;
   ( bdi_valid_bytes_3_port, bdi_valid_bytes_2_port, bdi_valid_bytes_1_port, 
      bdi_valid_bytes_0_port ) <= bdi_valid_bytes;
   ( bdi_size_2_port, bdi_size_1_port, bdi_size_0_port ) <= bdi_size;
   bdi_eot_port <= bdi_eot;
   decrypt_in_port <= decrypt_in;
   key_update_port <= key_update;
   hash_in_port <= hash_in;
   bdo <= ( bdo_31_port, bdo_30_port, bdo_29_port, bdo_28_port, bdo_27_port, 
      bdo_26_port, bdo_25_port, bdo_24_port, bdo_23_port, bdo_22_port, 
      bdo_21_port, bdo_20_port, bdo_19_port, bdo_18_port, bdo_17_port, 
      bdo_16_port, bdo_15_port, bdo_14_port, bdo_13_port, bdo_12_port, 
      bdo_11_port, bdo_10_port, bdo_9_port, bdo_8_port, bdo_7_port, bdo_6_port,
      bdo_5_port, bdo_4_port, bdo_3_port, bdo_2_port, bdo_1_port, bdo_0_port );
   bdo_valid <= bdo_valid_port;
   bdo_ready_port <= bdo_ready;
   bdo_type <= ( bdo_type_3_port, bdo_type_2_port, X_Logic0_port, bdo_type_0 );
   bdo_valid_bytes <= ( bdo_valid_bytes_3_port, bdo_valid_bytes_2_port, 
      bdo_valid_bytes_1_port, bdo_valid_bytes_0_port );
   end_of_block <= end_of_block_port;
   msg_auth_valid <= msg_auth_valid_port;
   msg_auth <= msg_auth_port;
   
   round_counter : counter_num_bits4_1 port map( clk => clk_port, reset => 
                           load_rnd, enable => en_rnd, q(3) => 
                           rnd_counter_3_port, q(2) => rnd_counter_2_port, q(1)
                           => rnd_counter_1_port, q(0) => rnd_counter_0_port);
   E_dcount : counter_num_bits4_1 port map( clk => clk_port, reset => 
                           load_dcount, enable => en_dcount, q(3) => 
                           dcount_3_port, q(2) => dcount_2_port, q(1) => 
                           dcount_1_port, q(0) => dcount_0_port);
   cyc_ops : cyclist_ops_DATA_LEN32_1 port map( clk => clk_port, key_en => 
                           key_en, state_main_en(2) => state_main_en_2_port, 
                           state_main_en(1) => state_main_en_1_port, 
                           state_main_en(0) => state_main_en_0_port, 
                           state_main_sel(6) => state_main_sel_6_port, 
                           state_main_sel(5) => state_main_sel_5_port, 
                           state_main_sel(4) => state_main_sel_4_port, 
                           state_main_sel(3) => state_main_sel_5_port, 
                           state_main_sel(2) => state_main_sel_2, 
                           state_main_sel(1) => state_main_sel_5_port, 
                           state_main_sel(0) => state_main_sel_0, 
                           cyc_state_update_sel => cyc_state_update_sel, 
                           xor_sel => xor_sel, cycd_sel(1) => cycd_sel_1_port, 
                           cycd_sel(0) => cycd_sel_0_port, extract_sel => 
                           extract_sel, bdi_key(31) => bdi_key_31_port, 
                           bdi_key(30) => bdi_key_30_port, bdi_key(29) => 
                           bdi_key_29_port, bdi_key(28) => bdi_key_28_port, 
                           bdi_key(27) => bdi_key_27_port, bdi_key(26) => 
                           bdi_key_26_port, bdi_key(25) => bdi_key_25_port, 
                           bdi_key(24) => bdi_key_24_port, bdi_key(23) => 
                           bdi_key_23_port, bdi_key(22) => bdi_key_22_port, 
                           bdi_key(21) => bdi_key_21_port, bdi_key(20) => 
                           bdi_key_20_port, bdi_key(19) => bdi_key_19_port, 
                           bdi_key(18) => bdi_key_18_port, bdi_key(17) => 
                           bdi_key_17_port, bdi_key(16) => bdi_key_16_port, 
                           bdi_key(15) => bdi_key_15_port, bdi_key(14) => 
                           bdi_key_14_port, bdi_key(13) => bdi_key_13_port, 
                           bdi_key(12) => bdi_key_12_port, bdi_key(11) => 
                           bdi_key_11_port, bdi_key(10) => bdi_key_10_port, 
                           bdi_key(9) => bdi_key_9_port, bdi_key(8) => 
                           bdi_key_8_port, bdi_key(7) => bdi_key_7_port, 
                           bdi_key(6) => bdi_key_6_port, bdi_key(5) => 
                           bdi_key_5_port, bdi_key(4) => bdi_key_4_port, 
                           bdi_key(3) => bdi_key_3_port, bdi_key(2) => 
                           bdi_key_2_port, bdi_key(1) => bdi_key_1_port, 
                           bdi_key(0) => bdi_key_0_port, cu_cd(7) => 
                           cu_cd_s_7_port, cu_cd(6) => cu_cd_s_6_port, cu_cd(5)
                           => X_Logic0_port, cu_cd(4) => X_Logic0_port, 
                           cu_cd(3) => X_Logic0_port, cu_cd(2) => X_Logic0_port
                           , cu_cd(1) => cu_cd_s_1, cu_cd(0) => cu_cd_s_0, 
                           dcount_in(3) => dcount_3_port, dcount_in(2) => 
                           dcount_2_port, dcount_in(1) => dcount_1_port, 
                           dcount_in(0) => dcount_0_port, rnd_counter(3) => 
                           rnd_counter_3_port, rnd_counter(2) => 
                           rnd_counter_2_port, rnd_counter(1) => 
                           rnd_counter_1_port, rnd_counter(0) => 
                           rnd_counter_0_port, bdo_out(31) => bdo_31_port, 
                           bdo_out(30) => bdo_30_port, bdo_out(29) => 
                           bdo_29_port, bdo_out(28) => bdo_28_port, bdo_out(27)
                           => bdo_27_port, bdo_out(26) => bdo_26_port, 
                           bdo_out(25) => bdo_25_port, bdo_out(24) => 
                           bdo_24_port, bdo_out(23) => bdo_23_port, bdo_out(22)
                           => bdo_22_port, bdo_out(21) => bdo_21_port, 
                           bdo_out(20) => bdo_20_port, bdo_out(19) => 
                           bdo_19_port, bdo_out(18) => bdo_18_port, bdo_out(17)
                           => bdo_17_port, bdo_out(16) => bdo_16_port, 
                           bdo_out(15) => bdo_15_port, bdo_out(14) => 
                           bdo_14_port, bdo_out(13) => bdo_13_port, bdo_out(12)
                           => bdo_12_port, bdo_out(11) => bdo_11_port, 
                           bdo_out(10) => bdo_10_port, bdo_out(9) => bdo_9_port
                           , bdo_out(8) => bdo_8_port, bdo_out(7) => bdo_7_port
                           , bdo_out(6) => bdo_6_port, bdo_out(5) => bdo_5_port
                           , bdo_out(4) => bdo_4_port, bdo_out(3) => bdo_3_port
                           , bdo_out(2) => bdo_2_port, bdo_out(1) => bdo_1_port
                           , bdo_out(0) => bdo_0_port);
   C30 : GTECH_AND2 port map( A => N76, B => N754, Z => N77);
   C31 : GTECH_AND2 port map( A => N77, B => N755, Z => N78);
   C33 : GTECH_OR2 port map( A => cyc_s_2_port, B => cyc_s_1_port, Z => N79);
   C34 : GTECH_OR2 port map( A => N79, B => N755, Z => N80);
   C37 : GTECH_OR2 port map( A => cyc_s_2_port, B => N754, Z => N82);
   C38 : GTECH_OR2 port map( A => N82, B => cyc_s_0_port, Z => N83);
   C42 : GTECH_OR2 port map( A => cyc_s_2_port, B => N754, Z => N85);
   C43 : GTECH_OR2 port map( A => N85, B => N755, Z => N86);
   C46 : GTECH_OR2 port map( A => N76, B => cyc_s_1_port, Z => N88);
   C47 : GTECH_OR2 port map( A => N88, B => cyc_s_0_port, Z => N89);
   C51 : GTECH_OR2 port map( A => N76, B => cyc_s_1_port, Z => N91);
   C52 : GTECH_OR2 port map( A => N91, B => N755, Z => N92);
   gt_294 : process ( X_Logic0_port, dcount_3_port, dcount_2_port, 
         dcount_1_port, dcount_0_port, X_Logic1_port )
      variable A : SIGNED( 31 downto 0 );
      variable B : SIGNED( 3 downto 0 );
      variable Z : SIGNED( 0 downto 0 );
   begin
      A := ( X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            dcount_3_port, dcount_2_port, dcount_1_port, dcount_0_port );
      B := ( X_Logic0_port, X_Logic1_port, X_Logic1_port, X_Logic1_port );
      if ( A > B ) then
         Z := ( others => '1' );
      else
         Z := ( others => '0' );
      end if;
      ( 0 => N196 ) <= Z;
   end process;
   
   gt_297 : process ( X_Logic0_port, dcount_3_port, dcount_2_port, 
         dcount_1_port, dcount_0_port, X_Logic1_port )
      variable A : SIGNED( 31 downto 0 );
      variable B : SIGNED( 2 downto 0 );
      variable Z : SIGNED( 0 downto 0 );
   begin
      A := ( X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            dcount_3_port, dcount_2_port, dcount_1_port, dcount_0_port );
      B := ( X_Logic0_port, X_Logic1_port, X_Logic1_port );
      if ( A > B ) then
         Z := ( others => '1' );
      else
         Z := ( others => '0' );
      end if;
      ( 0 => N198 ) <= Z;
   end process;
   
   gt_309 : process ( X_Logic0_port, dcount_3_port, dcount_2_port, 
         dcount_1_port, dcount_0_port, X_Logic1_port )
      variable A : SIGNED( 31 downto 0 );
      variable B : SIGNED( 3 downto 0 );
      variable Z : SIGNED( 0 downto 0 );
   begin
      A := ( X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            dcount_3_port, dcount_2_port, dcount_1_port, dcount_0_port );
      B := ( X_Logic0_port, X_Logic1_port, X_Logic1_port, X_Logic1_port );
      if ( A > B ) then
         Z := ( others => '1' );
      else
         Z := ( others => '0' );
      end if;
      ( 0 => N216 ) <= Z;
   end process;
   
   gt_312 : process ( X_Logic0_port, dcount_3_port, dcount_2_port, 
         dcount_1_port, dcount_0_port, X_Logic1_port )
      variable A : SIGNED( 31 downto 0 );
      variable B : SIGNED( 2 downto 0 );
      variable Z : SIGNED( 0 downto 0 );
   begin
      A := ( X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            dcount_3_port, dcount_2_port, dcount_1_port, dcount_0_port );
      B := ( X_Logic0_port, X_Logic1_port, X_Logic1_port );
      if ( A > B ) then
         Z := ( others => '1' );
      else
         Z := ( others => '0' );
      end if;
      ( 0 => N218 ) <= Z;
   end process;
   
   gt_341 : process ( X_Logic0_port, dcount_3_port, dcount_2_port, 
         dcount_1_port, dcount_0_port, X_Logic1_port )
      variable A : SIGNED( 31 downto 0 );
      variable B : SIGNED( 2 downto 0 );
      variable Z : SIGNED( 0 downto 0 );
   begin
      A := ( X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            dcount_3_port, dcount_2_port, dcount_1_port, dcount_0_port );
      B := ( X_Logic0_port, X_Logic1_port, X_Logic1_port );
      if ( A > B ) then
         Z := ( others => '1' );
      else
         Z := ( others => '0' );
      end if;
      ( 0 => N256 ) <= Z;
   end process;
   
   gt_355 : process ( X_Logic0_port, dcount_3_port, dcount_2_port, 
         dcount_1_port, dcount_0_port, X_Logic1_port )
      variable A : SIGNED( 31 downto 0 );
      variable B : SIGNED( 2 downto 0 );
      variable Z : SIGNED( 0 downto 0 );
   begin
      A := ( X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            dcount_3_port, dcount_2_port, dcount_1_port, dcount_0_port );
      B := ( X_Logic0_port, X_Logic1_port, X_Logic1_port );
      if ( A > B ) then
         Z := ( others => '1' );
      else
         Z := ( others => '0' );
      end if;
      ( 0 => N263 ) <= Z;
   end process;
   
   gt_382 : process ( X_Logic0_port, dcount_3_port, dcount_2_port, 
         dcount_1_port, dcount_0_port, X_Logic1_port )
      variable A : SIGNED( 31 downto 0 );
      variable B : SIGNED( 3 downto 0 );
      variable Z : SIGNED( 0 downto 0 );
   begin
      A := ( X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            dcount_3_port, dcount_2_port, dcount_1_port, dcount_0_port );
      B := ( X_Logic0_port, X_Logic1_port, X_Logic1_port, X_Logic1_port );
      if ( A > B ) then
         Z := ( others => '1' );
      else
         Z := ( others => '0' );
      end if;
      ( 0 => N323 ) <= Z;
   end process;
   
   gt_385 : process ( X_Logic0_port, dcount_3_port, dcount_2_port, 
         dcount_1_port, dcount_0_port, X_Logic1_port )
      variable A : SIGNED( 31 downto 0 );
      variable B : SIGNED( 2 downto 0 );
      variable Z : SIGNED( 0 downto 0 );
   begin
      A := ( X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            dcount_3_port, dcount_2_port, dcount_1_port, dcount_0_port );
      B := ( X_Logic0_port, X_Logic1_port, X_Logic1_port );
      if ( A > B ) then
         Z := ( others => '1' );
      else
         Z := ( others => '0' );
      end if;
      ( 0 => N325 ) <= Z;
   end process;
   
   lt_398 : process ( X_Logic0_port, dcount_3_port, dcount_2_port, 
         dcount_1_port, dcount_0_port, X_Logic1_port )
      variable A : SIGNED( 31 downto 0 );
      variable B : SIGNED( 4 downto 0 );
      variable Z : SIGNED( 0 downto 0 );
   begin
      A := ( X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            dcount_3_port, dcount_2_port, dcount_1_port, dcount_0_port );
      B := ( X_Logic0_port, X_Logic1_port, X_Logic0_port, X_Logic1_port, 
            X_Logic1_port );
      if ( A < B ) then
         Z := ( others => '1' );
      else
         Z := ( others => '0' );
      end if;
      ( 0 => N329 ) <= Z;
   end process;
   
   gt_421 : process ( X_Logic0_port, dcount_3_port, dcount_2_port, 
         dcount_1_port, dcount_0_port, X_Logic1_port )
      variable A : SIGNED( 31 downto 0 );
      variable B : SIGNED( 2 downto 0 );
      variable Z : SIGNED( 0 downto 0 );
   begin
      A := ( X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            dcount_3_port, dcount_2_port, dcount_1_port, dcount_0_port );
      B := ( X_Logic0_port, X_Logic1_port, X_Logic1_port );
      if ( A > B ) then
         Z := ( others => '1' );
      else
         Z := ( others => '0' );
      end if;
      ( 0 => N360 ) <= Z;
   end process;
   
   lt_426 : process ( X_Logic0_port, dcount_3_port, dcount_2_port, 
         dcount_1_port, dcount_0_port, X_Logic1_port )
      variable A : SIGNED( 31 downto 0 );
      variable B : SIGNED( 3 downto 0 );
      variable Z : SIGNED( 0 downto 0 );
   begin
      A := ( X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            dcount_3_port, dcount_2_port, dcount_1_port, dcount_0_port );
      B := ( X_Logic0_port, X_Logic1_port, X_Logic1_port, X_Logic0_port );
      if ( A < B ) then
         Z := ( others => '1' );
      else
         Z := ( others => '0' );
      end if;
      ( 0 => N363 ) <= Z;
   end process;
   
   gt_441 : process ( X_Logic0_port, dcount_3_port, dcount_2_port, 
         dcount_1_port, dcount_0_port, X_Logic1_port )
      variable A : SIGNED( 31 downto 0 );
      variable B : SIGNED( 2 downto 0 );
      variable Z : SIGNED( 0 downto 0 );
   begin
      A := ( X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            dcount_3_port, dcount_2_port, dcount_1_port, dcount_0_port );
      B := ( X_Logic0_port, X_Logic1_port, X_Logic1_port );
      if ( A > B ) then
         Z := ( others => '1' );
      else
         Z := ( others => '0' );
      end if;
      ( 0 => N369 ) <= Z;
   end process;
   
   gt_447 : process ( X_Logic0_port, dcount_3_port, dcount_2_port, 
         dcount_1_port, dcount_0_port, X_Logic1_port )
      variable A : SIGNED( 31 downto 0 );
      variable B : SIGNED( 2 downto 0 );
      variable Z : SIGNED( 0 downto 0 );
   begin
      A := ( X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            dcount_3_port, dcount_2_port, dcount_1_port, dcount_0_port );
      B := ( X_Logic0_port, X_Logic1_port, X_Logic1_port );
      if ( A > B ) then
         Z := ( others => '1' );
      else
         Z := ( others => '0' );
      end if;
      ( 0 => N371 ) <= Z;
   end process;
   
   ne_542 : process ( bdi_31_port, bdi_30_port, bdi_29_port, bdi_28_port, 
         bdi_27_port, bdi_26_port, bdi_25_port, bdi_24_port, bdi_23_port, 
         bdi_22_port, bdi_21_port, bdi_20_port, bdi_19_port, bdi_18_port, 
         bdi_17_port, bdi_16_port, bdi_15_port, bdi_14_port, bdi_13_port, 
         bdi_12_port, bdi_11_port, bdi_10_port, bdi_9_port, bdi_8_port, 
         bdi_7_port, bdi_6_port, bdi_5_port, bdi_4_port, bdi_3_port, bdi_2_port
         , bdi_1_port, bdi_0_port, bdo_31_port, bdo_30_port, bdo_29_port, 
         bdo_28_port, bdo_27_port, bdo_26_port, bdo_25_port, bdo_24_port, 
         bdo_23_port, bdo_22_port, bdo_21_port, bdo_20_port, bdo_19_port, 
         bdo_18_port, bdo_17_port, bdo_16_port, bdo_15_port, bdo_14_port, 
         bdo_13_port, bdo_12_port, bdo_11_port, bdo_10_port, bdo_9_port, 
         bdo_8_port, bdo_7_port, bdo_6_port, bdo_5_port, bdo_4_port, bdo_3_port
         , bdo_2_port, bdo_1_port, bdo_0_port )
      variable A : UNSIGNED( 31 downto 0 );
      variable B : UNSIGNED( 31 downto 0 );
      variable Z : UNSIGNED( 0 downto 0 );
   begin
      A := ( bdi_31_port, bdi_30_port, bdi_29_port, bdi_28_port, bdi_27_port, 
            bdi_26_port, bdi_25_port, bdi_24_port, bdi_23_port, bdi_22_port, 
            bdi_21_port, bdi_20_port, bdi_19_port, bdi_18_port, bdi_17_port, 
            bdi_16_port, bdi_15_port, bdi_14_port, bdi_13_port, bdi_12_port, 
            bdi_11_port, bdi_10_port, bdi_9_port, bdi_8_port, bdi_7_port, 
            bdi_6_port, bdi_5_port, bdi_4_port, bdi_3_port, bdi_2_port, 
            bdi_1_port, bdi_0_port );
      B := ( bdo_31_port, bdo_30_port, bdo_29_port, bdo_28_port, bdo_27_port, 
            bdo_26_port, bdo_25_port, bdo_24_port, bdo_23_port, bdo_22_port, 
            bdo_21_port, bdo_20_port, bdo_19_port, bdo_18_port, bdo_17_port, 
            bdo_16_port, bdo_15_port, bdo_14_port, bdo_13_port, bdo_12_port, 
            bdo_11_port, bdo_10_port, bdo_9_port, bdo_8_port, bdo_7_port, 
            bdo_6_port, bdo_5_port, bdo_4_port, bdo_3_port, bdo_2_port, 
            bdo_1_port, bdo_0_port );
      if ( A /= B ) then
         Z := ( others => '1' );
      else
         Z := ( others => '0' );
      end if;
      ( 0 => N546 ) <= Z;
   end process;
   
   ne_552 : process ( bdi_31_port, bdi_30_port, bdi_29_port, bdi_28_port, 
         bdi_27_port, bdi_26_port, bdi_25_port, bdi_24_port, bdi_23_port, 
         bdi_22_port, bdi_21_port, bdi_20_port, bdi_19_port, bdi_18_port, 
         bdi_17_port, bdi_16_port, bdi_15_port, bdi_14_port, bdi_13_port, 
         bdi_12_port, bdi_11_port, bdi_10_port, bdi_9_port, bdi_8_port, 
         bdi_7_port, bdi_6_port, bdi_5_port, bdi_4_port, bdi_3_port, bdi_2_port
         , bdi_1_port, bdi_0_port, bdo_31_port, bdo_30_port, bdo_29_port, 
         bdo_28_port, bdo_27_port, bdo_26_port, bdo_25_port, bdo_24_port, 
         bdo_23_port, bdo_22_port, bdo_21_port, bdo_20_port, bdo_19_port, 
         bdo_18_port, bdo_17_port, bdo_16_port, bdo_15_port, bdo_14_port, 
         bdo_13_port, bdo_12_port, bdo_11_port, bdo_10_port, bdo_9_port, 
         bdo_8_port, bdo_7_port, bdo_6_port, bdo_5_port, bdo_4_port, bdo_3_port
         , bdo_2_port, bdo_1_port, bdo_0_port )
      variable A : UNSIGNED( 31 downto 0 );
      variable B : UNSIGNED( 31 downto 0 );
      variable Z : UNSIGNED( 0 downto 0 );
   begin
      A := ( bdi_31_port, bdi_30_port, bdi_29_port, bdi_28_port, bdi_27_port, 
            bdi_26_port, bdi_25_port, bdi_24_port, bdi_23_port, bdi_22_port, 
            bdi_21_port, bdi_20_port, bdi_19_port, bdi_18_port, bdi_17_port, 
            bdi_16_port, bdi_15_port, bdi_14_port, bdi_13_port, bdi_12_port, 
            bdi_11_port, bdi_10_port, bdi_9_port, bdi_8_port, bdi_7_port, 
            bdi_6_port, bdi_5_port, bdi_4_port, bdi_3_port, bdi_2_port, 
            bdi_1_port, bdi_0_port );
      B := ( bdo_31_port, bdo_30_port, bdo_29_port, bdo_28_port, bdo_27_port, 
            bdo_26_port, bdo_25_port, bdo_24_port, bdo_23_port, bdo_22_port, 
            bdo_21_port, bdo_20_port, bdo_19_port, bdo_18_port, bdo_17_port, 
            bdo_16_port, bdo_15_port, bdo_14_port, bdo_13_port, bdo_12_port, 
            bdo_11_port, bdo_10_port, bdo_9_port, bdo_8_port, bdo_7_port, 
            bdo_6_port, bdo_5_port, bdo_4_port, bdo_3_port, bdo_2_port, 
            bdo_1_port, bdo_0_port );
      if ( A /= B ) then
         Z := ( others => '1' );
      else
         Z := ( others => '0' );
      end if;
      ( 0 => N549 ) <= Z;
   end process;
   
   bdi_eot_prev_reg : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => X_Logic1_port, next_state => N584
               , clocked_on => clk_port, Q => bdi_eot_prev, QN => n_1156);
   cyc_s_reg_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N594, next_state => N576, 
               clocked_on => clk_port, Q => cyc_s_2_port, QN => n_1157);
   cyc_s_reg_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N594, next_state => N575, 
               clocked_on => clk_port, Q => cyc_s_1_port, QN => n_1158);
   cyc_s_reg_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N594, next_state => N574, 
               clocked_on => clk_port, Q => cyc_s_0_port, QN => n_1159);
   mode_reg_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N603, next_state => X_Logic0_port
               , clocked_on => clk_port, Q => mode_1_port, QN => n_1160);
   mode_reg_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N603, next_state => N577, 
               clocked_on => clk_port, Q => mode_0_port, QN => n_1161);
   tag_verified_reg : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => X_Logic1_port, next_state => N578
               , clocked_on => clk_port, Q => tag_verified, QN => n_1162);
   calling_state_reg_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N611, next_state => N581, 
               clocked_on => clk_port, Q => calling_state_2_port, QN => n_1163
               );
   calling_state_reg_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N611, next_state => N580, 
               clocked_on => clk_port, Q => calling_state_1_port, QN => n_1164
               );
   calling_state_reg_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N611, next_state => N579, 
               clocked_on => clk_port, Q => calling_state_0_port, QN => n_1165
               );
   gtr_one_perm_reg : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N615, next_state => N582, 
               clocked_on => clk_port, Q => gtr_one_perm, QN => n_1166);
   decrypt_op_s_reg : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N621, next_state => N583, 
               clocked_on => clk_port, Q => decrypt_op_s, QN => n_1167);
   I_0 : GTECH_NOT port map( A => bdi_type(0), Z => N622);
   C1222 : GTECH_OR2 port map( A => N622, B => N638, Z => N623);
   I_1 : GTECH_NOT port map( A => N623, Z => N624);
   I_2 : GTECH_NOT port map( A => dcount_1_port, Z => N625);
   I_3 : GTECH_NOT port map( A => dcount_0_port, Z => N626);
   C1254 : GTECH_OR2 port map( A => dcount_2_port, B => dcount_3_port, Z => 
                           N627);
   C1255 : GTECH_OR2 port map( A => N625, B => N627, Z => N628);
   C1256 : GTECH_OR2 port map( A => N626, B => N628, Z => N629);
   I_4 : GTECH_NOT port map( A => N629, Z => N630);
   I_5 : GTECH_NOT port map( A => dcount_2_port, Z => N631);
   C1287 : GTECH_OR2 port map( A => N631, B => dcount_3_port, Z => N632);
   C1288 : GTECH_OR2 port map( A => dcount_1_port, B => N632, Z => N633);
   C1289 : GTECH_OR2 port map( A => dcount_0_port, B => N633, Z => N634);
   I_6 : GTECH_NOT port map( A => N634, Z => N635);
   I_7 : GTECH_NOT port map( A => bdi_type(2), Z => N636);
   C1292 : GTECH_OR2 port map( A => N636, B => bdi_type(3), Z => N637);
   C1293 : GTECH_OR2 port map( A => bdi_type(1), B => N637, Z => N638);
   C1294 : GTECH_OR2 port map( A => bdi_type(0), B => N638, Z => N639);
   I_8 : GTECH_NOT port map( A => N639, Z => N640);
   C1326 : GTECH_OR2 port map( A => dcount_2_port, B => dcount_3_port, Z => 
                           N641);
   C1327 : GTECH_OR2 port map( A => N625, B => N641, Z => N642);
   C1328 : GTECH_OR2 port map( A => N626, B => N642, Z => N643);
   I_9 : GTECH_NOT port map( A => N643, Z => N644);
   I_10 : GTECH_NOT port map( A => calling_state_2_port, Z => N645);
   I_11 : GTECH_NOT port map( A => calling_state_1_port, Z => N646);
   C1332 : GTECH_OR2 port map( A => N646, B => N645, Z => N647);
   C1333 : GTECH_OR2 port map( A => calling_state_0_port, B => N647, Z => N648)
                           ;
   I_12 : GTECH_NOT port map( A => N648, Z => N649);
   I_13 : GTECH_NOT port map( A => mode_0_port, Z => N650);
   C1336 : GTECH_OR2 port map( A => N650, B => mode_1_port, Z => N651);
   I_14 : GTECH_NOT port map( A => N651, Z => N652);
   C1339 : GTECH_OR2 port map( A => calling_state_1_port, B => N645, Z => N653)
                           ;
   C1340 : GTECH_OR2 port map( A => calling_state_0_port, B => N653, Z => N654)
                           ;
   C1343 : GTECH_AND2 port map( A => bdi_valid_bytes_2_port, B => 
                           bdi_valid_bytes_3_port, Z => N655);
   C1344 : GTECH_AND2 port map( A => bdi_valid_bytes_1_port, B => N655, Z => 
                           N656);
   C1345 : GTECH_AND2 port map( A => bdi_valid_bytes_0_port, B => N656, Z => 
                           N657);
   I_15 : GTECH_NOT port map( A => bdi_size_2_port, Z => N658);
   C1347 : GTECH_OR2 port map( A => bdi_size_1_port, B => N658, Z => N659);
   C1348 : GTECH_OR2 port map( A => bdi_size_0_port, B => N659, Z => N660);
   I_16 : GTECH_NOT port map( A => N660, Z => N661);
   C1380 : GTECH_OR2 port map( A => dcount_2_port, B => dcount_3_port, Z => 
                           N662);
   C1381 : GTECH_OR2 port map( A => N625, B => N662, Z => N663);
   C1382 : GTECH_OR2 port map( A => N626, B => N663, Z => N664);
   I_17 : GTECH_NOT port map( A => N664, Z => N665);
   I_18 : GTECH_NOT port map( A => dcount_3_port, Z => N666);
   C1415 : GTECH_OR2 port map( A => dcount_2_port, B => N666, Z => N667);
   C1416 : GTECH_OR2 port map( A => N625, B => N667, Z => N668);
   C1417 : GTECH_OR2 port map( A => N626, B => N668, Z => N669);
   I_19 : GTECH_NOT port map( A => N669, Z => N670);
   C1456 : GTECH_OR2 port map( A => N631, B => dcount_3_port, Z => N671);
   C1457 : GTECH_OR2 port map( A => dcount_1_port, B => N671, Z => N672);
   C1458 : GTECH_OR2 port map( A => N626, B => N672, Z => N673);
   I_20 : GTECH_NOT port map( A => N673, Z => N674);
   C1497 : GTECH_OR2 port map( A => dcount_2_port, B => dcount_3_port, Z => 
                           N675);
   C1498 : GTECH_OR2 port map( A => N625, B => N675, Z => N676);
   C1499 : GTECH_OR2 port map( A => N626, B => N676, Z => N677);
   I_21 : GTECH_NOT port map( A => N677, Z => N678);
   C1531 : GTECH_OR2 port map( A => dcount_2_port, B => dcount_3_port, Z => 
                           N679);
   C1532 : GTECH_OR2 port map( A => N625, B => N679, Z => N680);
   C1533 : GTECH_OR2 port map( A => N626, B => N680, Z => N681);
   I_22 : GTECH_NOT port map( A => N681, Z => N682);
   I_23 : GTECH_NOT port map( A => calling_state_0_port, Z => N683);
   C1537 : GTECH_OR2 port map( A => N646, B => calling_state_2_port, Z => N684)
                           ;
   C1538 : GTECH_OR2 port map( A => N683, B => N684, Z => N685);
   I_24 : GTECH_NOT port map( A => N685, Z => N686);
   C1541 : GTECH_OR2 port map( A => calling_state_1_port, B => N645, Z => N687)
                           ;
   C1542 : GTECH_OR2 port map( A => calling_state_0_port, B => N687, Z => N688)
                           ;
   I_25 : GTECH_NOT port map( A => N688, Z => N689);
   C1573 : GTECH_OR2 port map( A => N631, B => dcount_3_port, Z => N690);
   C1574 : GTECH_OR2 port map( A => dcount_1_port, B => N690, Z => N691);
   C1575 : GTECH_OR2 port map( A => dcount_0_port, B => N691, Z => N692);
   C1613 : GTECH_OR2 port map( A => dcount_2_port, B => dcount_3_port, Z => 
                           N693);
   C1614 : GTECH_OR2 port map( A => N625, B => N693, Z => N694);
   C1615 : GTECH_OR2 port map( A => N626, B => N694, Z => N695);
   I_26 : GTECH_NOT port map( A => N695, Z => N696);
   C1619 : GTECH_OR2 port map( A => calling_state_1_port, B => N645, Z => N697)
                           ;
   C1620 : GTECH_OR2 port map( A => N683, B => N697, Z => N698);
   I_27 : GTECH_NOT port map( A => N698, Z => N699);
   I_28 : GTECH_NOT port map( A => rnd_counter_3_port, Z => N700);
   I_29 : GTECH_NOT port map( A => rnd_counter_1_port, Z => N701);
   I_30 : GTECH_NOT port map( A => rnd_counter_0_port, Z => N702);
   C1625 : GTECH_OR2 port map( A => rnd_counter_2_port, B => N700, Z => N703);
   C1626 : GTECH_OR2 port map( A => N701, B => N703, Z => N704);
   C1627 : GTECH_OR2 port map( A => N702, B => N704, Z => N705);
   I_31 : GTECH_NOT port map( A => N705, Z => N706);
   C1629 : GTECH_OR2 port map( A => bdi_size_0_port, B => bdi_size_1_port, Z =>
                           N707);
   I_32 : GTECH_NOT port map( A => decrypt_op_s, Z => N708);
   C1688 : GTECH_OR2 port map( A => dcount_2_port, B => N666, Z => N709);
   C1689 : GTECH_OR2 port map( A => N625, B => N709, Z => N710);
   C1690 : GTECH_OR2 port map( A => dcount_0_port, B => N710, Z => N711);
   I_33 : GTECH_NOT port map( A => N711, Z => N712);
   C1693 : GTECH_OR2 port map( A => calling_state_1_port, B => 
                           calling_state_2_port, Z => N713);
   C1694 : GTECH_OR2 port map( A => N683, B => N713, Z => N714);
   I_34 : GTECH_NOT port map( A => N714, Z => N715);
   C1698 : GTECH_OR2 port map( A => calling_state_1_port, B => N645, Z => N716)
                           ;
   C1699 : GTECH_OR2 port map( A => N683, B => N716, Z => N717);
   I_35 : GTECH_NOT port map( A => N717, Z => N718);
   C1721 : GTECH_OR2 port map( A => bdi_type(2), B => bdi_type(3), Z => N719);
   C1722 : GTECH_OR2 port map( A => bdi_type(1), B => N719, Z => N720);
   C1723 : GTECH_OR2 port map( A => N622, B => N720, Z => N721);
   I_36 : GTECH_NOT port map( A => N721, Z => N722);
   C1727 : GTECH_OR2 port map( A => bdi_type(0), B => N720, Z => N723);
   I_37 : GTECH_NOT port map( A => N723, Z => N724);
   I_38 : GTECH_NOT port map( A => bdi_type(1), Z => N725);
   C1733 : GTECH_OR2 port map( A => N725, B => N637, Z => N726);
   C1734 : GTECH_OR2 port map( A => N622, B => N726, Z => N727);
   I_39 : GTECH_NOT port map( A => N727, Z => N728);
   C1737 : GTECH_OR2 port map( A => N646, B => calling_state_2_port, Z => N729)
                           ;
   C1738 : GTECH_OR2 port map( A => calling_state_0_port, B => N729, Z => N730)
                           ;
   I_40 : GTECH_NOT port map( A => N730, Z => N731);
   C1741 : GTECH_OR2 port map( A => calling_state_1_port, B => 
                           calling_state_2_port, Z => N732);
   C1742 : GTECH_OR2 port map( A => N683, B => N732, Z => N733);
   I_41 : GTECH_NOT port map( A => N733, Z => N734);
   C1746 : GTECH_OR2 port map( A => calling_state_1_port, B => N645, Z => N735)
                           ;
   C1747 : GTECH_OR2 port map( A => N683, B => N735, Z => N736);
   I_42 : GTECH_NOT port map( A => N736, Z => N737);
   C1750 : GTECH_OR2 port map( A => calling_state_1_port, B => 
                           calling_state_2_port, Z => N738);
   C1751 : GTECH_OR2 port map( A => N683, B => N738, Z => N739);
   I_43 : GTECH_NOT port map( A => N739, Z => N740);
   C1753 : GTECH_OR2 port map( A => calling_state_1_port, B => 
                           calling_state_2_port, Z => N741);
   C1754 : GTECH_OR2 port map( A => calling_state_0_port, B => N741, Z => N742)
                           ;
   I_44 : GTECH_NOT port map( A => N742, Z => N743);
   C1756 : GTECH_OR2 port map( A => bdi_valid_bytes_2_port, B => 
                           bdi_valid_bytes_3_port, Z => N744);
   C1757 : GTECH_OR2 port map( A => bdi_valid_bytes_1_port, B => N744, Z => 
                           N745);
   C1758 : GTECH_OR2 port map( A => bdi_valid_bytes_0_port, B => N745, Z => 
                           N746);
   I_45 : GTECH_NOT port map( A => N746, Z => N747);
   C1760 : GTECH_OR2 port map( A => calling_state_1_port, B => 
                           calling_state_2_port, Z => N748);
   C1761 : GTECH_OR2 port map( A => calling_state_0_port, B => N748, Z => N749)
                           ;
   I_46 : GTECH_NOT port map( A => N749, Z => N750);
   I_47 : GTECH_NOT port map( A => bdi_eot_prev, Z => N751);
   I_48 : GTECH_NOT port map( A => bdi_eot_port, Z => N752);
   I_49 : GTECH_NOT port map( A => gtr_one_perm, Z => N753);
   I_50 : GTECH_NOT port map( A => cyc_s_1_port, Z => N754);
   I_51 : GTECH_NOT port map( A => cyc_s_0_port, Z => N755);
   C1784 : GTECH_OR2 port map( A => N754, B => cyc_s_2_port, Z => N756);
   C1785 : GTECH_OR2 port map( A => N755, B => N756, Z => N757);
   I_52 : GTECH_NOT port map( A => N757, Z => N758);
   C1801 : GTECH_OR2 port map( A => X_Logic0_port, B => X_Logic0_port, Z => 
                           N759);
   C1802 : GTECH_OR2 port map( A => X_Logic0_port, B => N759, Z => N760);
   C1803 : GTECH_OR2 port map( A => X_Logic0_port, B => N760, Z => N761);
   C1804 : GTECH_OR2 port map( A => X_Logic0_port, B => N761, Z => N762);
   C1805 : GTECH_OR2 port map( A => X_Logic0_port, B => N762, Z => N763);
   C1806 : GTECH_OR2 port map( A => X_Logic0_port, B => N763, Z => N764);
   C1807 : GTECH_OR2 port map( A => X_Logic0_port, B => N764, Z => N765);
   C1808 : GTECH_OR2 port map( A => X_Logic0_port, B => N765, Z => N766);
   C1809 : GTECH_OR2 port map( A => X_Logic0_port, B => N766, Z => N767);
   C1810 : GTECH_OR2 port map( A => X_Logic0_port, B => N767, Z => N768);
   C1811 : GTECH_OR2 port map( A => X_Logic0_port, B => N768, Z => N769);
   C1812 : GTECH_OR2 port map( A => X_Logic0_port, B => N769, Z => N770);
   C1813 : GTECH_OR2 port map( A => X_Logic0_port, B => N770, Z => N771);
   C1814 : GTECH_OR2 port map( A => X_Logic0_port, B => N771, Z => N772);
   C1815 : GTECH_OR2 port map( A => X_Logic0_port, B => N772, Z => N773);
   C1816 : GTECH_OR2 port map( A => X_Logic0_port, B => N773, Z => N774);
   C1817 : GTECH_OR2 port map( A => X_Logic0_port, B => N774, Z => N775);
   C1818 : GTECH_OR2 port map( A => X_Logic0_port, B => N775, Z => N776);
   C1819 : GTECH_OR2 port map( A => X_Logic0_port, B => N776, Z => N777);
   C1820 : GTECH_OR2 port map( A => X_Logic0_port, B => N777, Z => N778);
   C1821 : GTECH_OR2 port map( A => X_Logic0_port, B => N778, Z => N779);
   C1822 : GTECH_OR2 port map( A => X_Logic0_port, B => N779, Z => N780);
   C1823 : GTECH_OR2 port map( A => X_Logic0_port, B => N780, Z => N781);
   C1824 : GTECH_OR2 port map( A => X_Logic0_port, B => N781, Z => N782);
   C1825 : GTECH_OR2 port map( A => X_Logic0_port, B => N782, Z => N783);
   C1826 : GTECH_OR2 port map( A => X_Logic0_port, B => N783, Z => N784);
   C1827 : GTECH_OR2 port map( A => X_Logic0_port, B => N784, Z => N785);
   C1828 : GTECH_OR2 port map( A => dcount_3_port, B => N785, Z => N786);
   C1829 : GTECH_OR2 port map( A => N631, B => N786, Z => N787);
   C1830 : GTECH_OR2 port map( A => N625, B => N787, Z => N788);
   C1831 : GTECH_OR2 port map( A => dcount_0_port, B => N788, Z => N789);
   I_53 : GTECH_NOT port map( A => N789, Z => N790);
   C1861 : GTECH_OR2 port map( A => dcount_3_port, B => N785, Z => N791);
   C1862 : GTECH_OR2 port map( A => N631, B => N791, Z => N792);
   C1863 : GTECH_OR2 port map( A => dcount_1_port, B => N792, Z => N793);
   C1864 : GTECH_OR2 port map( A => dcount_0_port, B => N793, Z => N794);
   C1895 : GTECH_OR2 port map( A => dcount_3_port, B => N785, Z => N795);
   C1896 : GTECH_OR2 port map( A => N631, B => N795, Z => N796);
   C1897 : GTECH_OR2 port map( A => dcount_1_port, B => N796, Z => N797);
   C1898 : GTECH_OR2 port map( A => dcount_0_port, B => N797, Z => N798);
   C1902 : GTECH_OR2 port map( A => calling_state_1_port, B => N645, Z => N799)
                           ;
   C1903 : GTECH_OR2 port map( A => calling_state_0_port, B => N799, Z => N800)
                           ;
   I_54 : GTECH_NOT port map( A => N800, Z => N801);
   C1906_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic1_port, 
         -- Connections to port 'DATA2'
         DATA(1) => N624, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N0, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N1, 
         -- Connections to port 'Z'
         Z(0) => extract_sel );
   B_0 : GTECH_BUF port map( A => N640, Z => N0);
   B_1 : GTECH_BUF port map( A => N639, Z => N1);
   C1907_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 3 )
      port map(
         -- Connections to port 'DATA1'
         DATA(2) => X_Logic0_port, DATA(1) => X_Logic1_port, DATA(0) => 
               X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(5) => N623, DATA(4) => N624, DATA(3) => N624, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N0, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N1, 
         -- Connections to port 'Z'
         Z(2) => bdo_type_3_port, Z(1) => bdo_type_2_port, Z(0) => bdo_type_0 
               );
   C1908_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 2 )
      port map(
         -- Connections to port 'DATA1'
         DATA(1) => X_Logic1_port, DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(3) => N97, DATA(2) => key_update_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N2, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N3, 
         -- Connections to port 'Z'
         Z(1) => N99, Z(0) => N98 );
   B_2 : GTECH_BUF port map( A => hash_in_port, Z => N2);
   B_3 : GTECH_BUF port map( A => N96, Z => N3);
   C1909_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic1_port, 
         -- Connections to port 'DATA2'
         DATA(1) => key_update_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N2, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N3, 
         -- Connections to port 'Z'
         Z(0) => N100 );
   C1910_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => N100, 
         -- Connections to port 'DATA2'
         DATA(1) => X_Logic1_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N4, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N95, 
         -- Connections to port 'Z'
         Z(0) => N101 );
   B_4 : GTECH_BUF port map( A => N94, Z => N4);
   C1911_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 32 )
      port map(
         -- Connections to port 'DATA1'
         DATA(31) => X_Logic0_port, DATA(30) => X_Logic0_port, DATA(29) => 
               X_Logic0_port, DATA(28) => X_Logic0_port, DATA(27) => 
               X_Logic0_port, DATA(26) => X_Logic0_port, DATA(25) => 
               X_Logic0_port, DATA(24) => X_Logic0_port, DATA(23) => 
               X_Logic0_port, DATA(22) => X_Logic0_port, DATA(21) => 
               X_Logic0_port, DATA(20) => X_Logic0_port, DATA(19) => 
               X_Logic0_port, DATA(18) => X_Logic0_port, DATA(17) => 
               X_Logic0_port, DATA(16) => X_Logic1_port, DATA(15) => 
               X_Logic0_port, DATA(14) => X_Logic0_port, DATA(13) => 
               X_Logic0_port, DATA(12) => X_Logic0_port, DATA(11) => 
               X_Logic0_port, DATA(10) => X_Logic0_port, DATA(9) => 
               X_Logic0_port, DATA(8) => X_Logic0_port, DATA(7) => 
               X_Logic0_port, DATA(6) => X_Logic0_port, DATA(5) => 
               X_Logic0_port, DATA(4) => X_Logic0_port, DATA(3) => 
               X_Logic0_port, DATA(2) => X_Logic0_port, DATA(1) => 
               X_Logic0_port, DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(63) => bdi_31_port, DATA(62) => bdi_30_port, DATA(61) => 
               bdi_29_port, DATA(60) => bdi_28_port, DATA(59) => bdi_27_port, 
               DATA(58) => bdi_26_port, DATA(57) => bdi_25_port, DATA(56) => 
               bdi_24_port, DATA(55) => bdi_23_port, DATA(54) => bdi_22_port, 
               DATA(53) => bdi_21_port, DATA(52) => bdi_20_port, DATA(51) => 
               bdi_19_port, DATA(50) => bdi_18_port, DATA(49) => bdi_17_port, 
               DATA(48) => bdi_16_port, DATA(47) => bdi_15_port, DATA(46) => 
               bdi_14_port, DATA(45) => bdi_13_port, DATA(44) => bdi_12_port, 
               DATA(43) => bdi_11_port, DATA(42) => bdi_10_port, DATA(41) => 
               bdi_9_port, DATA(40) => bdi_8_port, DATA(39) => bdi_7_port, 
               DATA(38) => bdi_6_port, DATA(37) => bdi_5_port, DATA(36) => 
               bdi_4_port, DATA(35) => bdi_3_port, DATA(34) => bdi_2_port, 
               DATA(33) => bdi_1_port, DATA(32) => bdi_0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N5, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N6, 
         -- Connections to port 'Z'
         Z(31) => N134, Z(30) => N133, Z(29) => N132, Z(28) => N131, Z(27) => 
               N130, Z(26) => N129, Z(25) => N128, Z(24) => N127, Z(23) => N126
               , Z(22) => N125, Z(21) => N124, Z(20) => N123, Z(19) => N122, 
               Z(18) => N121, Z(17) => N120, Z(16) => N119, Z(15) => N118, 
               Z(14) => N117, Z(13) => N116, Z(12) => N115, Z(11) => N114, 
               Z(10) => N113, Z(9) => N112, Z(8) => N111, Z(7) => N110, Z(6) =>
               N109, Z(5) => N108, Z(4) => N107, Z(3) => N106, Z(2) => N105, 
               Z(1) => N104, Z(0) => N103 );
   B_5 : GTECH_BUF port map( A => N635, Z => N5);
   B_6 : GTECH_BUF port map( A => N634, Z => N6);
   C1912_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 3 )
      port map(
         -- Connections to port 'DATA1'
         DATA(2) => X_Logic1_port, DATA(1) => X_Logic0_port, DATA(0) => 
               X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(5) => cyc_s_2_port, DATA(4) => cyc_s_1_port, DATA(3) => 
               cyc_s_0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N5, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N6, 
         -- Connections to port 'Z'
         Z(2) => N137, Z(1) => N136, Z(0) => N135 );
   C1913_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 3 )
      port map(
         -- Connections to port 'DATA1'
         DATA(2) => X_Logic1_port, DATA(1) => X_Logic1_port, DATA(0) => 
               X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(5) => calling_state_2_port, DATA(4) => calling_state_1_port, 
               DATA(3) => calling_state_0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N5, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N6, 
         -- Connections to port 'Z'
         Z(2) => N140, Z(1) => N139, Z(0) => N138 );
   C1914_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 32 )
      port map(
         -- Connections to port 'DATA1'
         DATA(31) => key_31_port, DATA(30) => key_30_port, DATA(29) => 
               key_29_port, DATA(28) => key_28_port, DATA(27) => key_27_port, 
               DATA(26) => key_26_port, DATA(25) => key_25_port, DATA(24) => 
               key_24_port, DATA(23) => key_23_port, DATA(22) => key_22_port, 
               DATA(21) => key_21_port, DATA(20) => key_20_port, DATA(19) => 
               key_19_port, DATA(18) => key_18_port, DATA(17) => key_17_port, 
               DATA(16) => key_16_port, DATA(15) => key_15_port, DATA(14) => 
               key_14_port, DATA(13) => key_13_port, DATA(12) => key_12_port, 
               DATA(11) => key_11_port, DATA(10) => key_10_port, DATA(9) => 
               key_9_port, DATA(8) => key_8_port, DATA(7) => key_7_port, 
               DATA(6) => key_6_port, DATA(5) => key_5_port, DATA(4) => 
               key_4_port, DATA(3) => key_3_port, DATA(2) => key_2_port, 
               DATA(1) => key_1_port, DATA(0) => key_0_port, 
         -- Connections to port 'DATA2'
         DATA(63) => N134, DATA(62) => N133, DATA(61) => N132, DATA(60) => N131
               , DATA(59) => N130, DATA(58) => N129, DATA(57) => N128, DATA(56)
               => N127, DATA(55) => N126, DATA(54) => N125, DATA(53) => N124, 
               DATA(52) => N123, DATA(51) => N122, DATA(50) => N121, DATA(49) 
               => N120, DATA(48) => N119, DATA(47) => N118, DATA(46) => N117, 
               DATA(45) => N116, DATA(44) => N115, DATA(43) => N114, DATA(42) 
               => N113, DATA(41) => N112, DATA(40) => N111, DATA(39) => N110, 
               DATA(38) => N109, DATA(37) => N108, DATA(36) => N107, DATA(35) 
               => N106, DATA(34) => N105, DATA(33) => N104, DATA(32) => N103, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N7, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N8, 
         -- Connections to port 'Z'
         Z(31) => N172, Z(30) => N171, Z(29) => N170, Z(28) => N169, Z(27) => 
               N168, Z(26) => N167, Z(25) => N166, Z(24) => N165, Z(23) => N164
               , Z(22) => N163, Z(21) => N162, Z(20) => N161, Z(19) => N160, 
               Z(18) => N159, Z(17) => N158, Z(16) => N157, Z(15) => N156, 
               Z(14) => N155, Z(13) => N154, Z(12) => N153, Z(11) => N152, 
               Z(10) => N151, Z(9) => N150, Z(8) => N149, Z(7) => N148, Z(6) =>
               N147, Z(5) => N146, Z(4) => N145, Z(3) => N144, Z(2) => N143, 
               Z(1) => N142, Z(0) => N141 );
   B_7 : GTECH_BUF port map( A => key_valid_port, Z => N7);
   B_8 : GTECH_BUF port map( A => N102, Z => N8);
   C1915_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => N635, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N7, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N8, 
         -- Connections to port 'Z'
         Z(0) => N173 );
   C1916_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 3 )
      port map(
         -- Connections to port 'DATA1'
         DATA(2) => X_Logic0_port, DATA(1) => X_Logic1_port, DATA(0) => 
               X_Logic1_port, 
         -- Connections to port 'DATA2'
         DATA(5) => cyc_s_2_port, DATA(4) => cyc_s_1_port, DATA(3) => 
               cyc_s_0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N9, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N10, 
         -- Connections to port 'Z'
         Z(2) => N178, Z(1) => N177, Z(0) => N176 );
   B_9 : GTECH_BUF port map( A => N644, Z => N9);
   B_10 : GTECH_BUF port map( A => N643, Z => N10);
   C1917_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 3 )
      port map(
         -- Connections to port 'DATA1'
         DATA(2) => N178, DATA(1) => N177, DATA(0) => N176, 
         -- Connections to port 'DATA2'
         DATA(5) => cyc_s_2_port, DATA(4) => cyc_s_1_port, DATA(3) => 
               cyc_s_0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N11, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N12, 
         -- Connections to port 'Z'
         Z(2) => N181, Z(1) => N180, Z(0) => N179 );
   B_11 : GTECH_BUF port map( A => bdi_valid_port, Z => N11);
   B_12 : GTECH_BUF port map( A => N175, Z => N12);
   I_55 : GTECH_NOT port map( A => N198, Z => N199);
   C1919_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 2 )
      port map(
         -- Connections to port 'DATA1'
         DATA(1) => X_Logic0_port, DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(3) => N198, DATA(2) => N199, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N13, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N197, 
         -- Connections to port 'Z'
         Z(1) => N201, Z(0) => N200 );
   B_13 : GTECH_BUF port map( A => N196, Z => N13);
   C1920_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 2 )
      port map(
         -- Connections to port 'DATA1'
         DATA(1) => N201, DATA(0) => N200, 
         -- Connections to port 'DATA2'
         DATA(3) => X_Logic0_port, DATA(2) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N14, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N194, 
         -- Connections to port 'Z'
         Z(1) => N203, Z(0) => N202 );
   B_14 : GTECH_BUF port map( A => N657, Z => N14);
   C1921_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => N196, 
         -- Connections to port 'DATA2'
         DATA(1) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N14, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N194, 
         -- Connections to port 'Z'
         Z(0) => N204 );
   C1922_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 3 )
      port map(
         -- Connections to port 'DATA1'
         DATA(2) => X_Logic0_port, DATA(1) => X_Logic1_port, DATA(0) => 
               X_Logic1_port, 
         -- Connections to port 'DATA2'
         DATA(5) => cyc_s_2_port, DATA(4) => cyc_s_1_port, DATA(3) => 
               cyc_s_0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N15, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N209, 
         -- Connections to port 'Z'
         Z(2) => N212, Z(1) => N211, Z(0) => N210 );
   B_15 : GTECH_BUF port map( A => N208, Z => N15);
   C1923_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 3 )
      port map(
         -- Connections to port 'DATA1'
         DATA(2) => X_Logic0_port, DATA(1) => X_Logic1_port, DATA(0) => 
               X_Logic1_port, 
         -- Connections to port 'DATA2'
         DATA(5) => N212, DATA(4) => N211, DATA(3) => N210, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N16, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N207, 
         -- Connections to port 'Z'
         Z(2) => N215, Z(1) => N214, Z(0) => N213 );
   B_16 : GTECH_BUF port map( A => N206, Z => N16);
   I_56 : GTECH_NOT port map( A => N218, Z => N219);
   C1925_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 2 )
      port map(
         -- Connections to port 'DATA1'
         DATA(1) => X_Logic0_port, DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(3) => N218, DATA(2) => N219, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N17, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N217, 
         -- Connections to port 'Z'
         Z(1) => N221, Z(0) => N220 );
   B_17 : GTECH_BUF port map( A => N216, Z => N17);
   C1926_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 3 )
      port map(
         -- Connections to port 'DATA1'
         DATA(2) => X_Logic0_port, DATA(1) => X_Logic1_port, DATA(0) => 
               X_Logic1_port, 
         -- Connections to port 'DATA2'
         DATA(5) => N215, DATA(4) => N214, DATA(3) => N213, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N18, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N19, 
         -- Connections to port 'Z'
         Z(2) => N224, Z(1) => N223, Z(0) => N222 );
   B_18 : GTECH_BUF port map( A => bdi_eot_port, Z => N18);
   B_19 : GTECH_BUF port map( A => N752, Z => N19);
   C1927_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => N204, 
         -- Connections to port 'DATA2'
         DATA(1) => N216, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N18, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N19, 
         -- Connections to port 'Z'
         Z(0) => N225 );
   C1928_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => N657, 
         -- Connections to port 'DATA2'
         DATA(1) => X_Logic1_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N18, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N19, 
         -- Connections to port 'Z'
         Z(0) => N226 );
   C1929_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 2 )
      port map(
         -- Connections to port 'DATA1'
         DATA(1) => N203, DATA(0) => N202, 
         -- Connections to port 'DATA2'
         DATA(3) => N221, DATA(2) => N220, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N18, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N19, 
         -- Connections to port 'Z'
         Z(1) => N228, Z(0) => N227 );
   C1930_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 3 )
      port map(
         -- Connections to port 'DATA1'
         DATA(2) => X_Logic0_port, DATA(1) => X_Logic1_port, DATA(0) => 
               X_Logic1_port, 
         -- Connections to port 'DATA2'
         DATA(5) => cyc_s_2_port, DATA(4) => cyc_s_1_port, DATA(3) => 
               cyc_s_0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N20, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N230, 
         -- Connections to port 'Z'
         Z(2) => N233, Z(1) => N232, Z(0) => N231 );
   B_20 : GTECH_BUF port map( A => N229, Z => N20);
   C1931_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 2 )
      port map(
         -- Connections to port 'DATA1'
         DATA(1) => N228, DATA(0) => N227, 
         -- Connections to port 'DATA2'
         DATA(3) => X_Logic0_port, DATA(2) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N11, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N12, 
         -- Connections to port 'Z'
         Z(1) => N235, Z(0) => N234 );
   C1932_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 3 )
      port map(
         -- Connections to port 'DATA1'
         DATA(2) => N224, DATA(1) => N223, DATA(0) => N222, 
         -- Connections to port 'DATA2'
         DATA(5) => N233, DATA(4) => N232, DATA(3) => N231, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N11, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N12, 
         -- Connections to port 'Z'
         Z(2) => N238, Z(1) => N237, Z(0) => N236 );
   C1933_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => N225, 
         -- Connections to port 'DATA2'
         DATA(1) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N11, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N12, 
         -- Connections to port 'Z'
         Z(0) => N239 );
   C1934_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => N226, 
         -- Connections to port 'DATA2'
         DATA(1) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N11, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N12, 
         -- Connections to port 'Z'
         Z(0) => N240 );
   C1935_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => N240, 
         -- Connections to port 'DATA2'
         DATA(1) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N21, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N190, 
         -- Connections to port 'Z'
         Z(0) => N241 );
   B_21 : GTECH_BUF port map( A => N189, Z => N21);
   C1936_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 2 )
      port map(
         -- Connections to port 'DATA1'
         DATA(1) => N235, DATA(0) => N234, 
         -- Connections to port 'DATA2'
         DATA(3) => X_Logic0_port, DATA(2) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N21, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N190, 
         -- Connections to port 'Z'
         Z(1) => N243, Z(0) => N242 );
   C1937_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 3 )
      port map(
         -- Connections to port 'DATA1'
         DATA(2) => N238, DATA(1) => N237, DATA(0) => N236, 
         -- Connections to port 'DATA2'
         DATA(5) => X_Logic0_port, DATA(4) => X_Logic1_port, DATA(3) => 
               X_Logic1_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N21, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N190, 
         -- Connections to port 'Z'
         Z(2) => N246, Z(1) => N245, Z(0) => N244 );
   C1938_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => N239, 
         -- Connections to port 'DATA2'
         DATA(1) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N21, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N190, 
         -- Connections to port 'Z'
         Z(0) => N247 );
   I_57 : GTECH_NOT port map( A => N256, Z => N257);
   C1940_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 2 )
      port map(
         -- Connections to port 'DATA1'
         DATA(1) => N256, DATA(0) => N257, 
         -- Connections to port 'DATA2'
         DATA(3) => X_Logic0_port, DATA(2) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N22, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N23, 
         -- Connections to port 'Z'
         Z(1) => N259, Z(0) => N258 );
   B_22 : GTECH_BUF port map( A => N661, Z => N22);
   B_23 : GTECH_BUF port map( A => N660, Z => N23);
   C1941_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 3 )
      port map(
         -- Connections to port 'DATA1'
         DATA(2) => X_Logic0_port, DATA(1) => X_Logic1_port, DATA(0) => 
               X_Logic1_port, 
         -- Connections to port 'DATA2'
         DATA(5) => cyc_s_2_port, DATA(4) => cyc_s_1_port, DATA(3) => 
               cyc_s_0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N24, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N25, 
         -- Connections to port 'Z'
         Z(2) => N262, Z(1) => N261, Z(0) => N260 );
   B_24 : GTECH_BUF port map( A => N674, Z => N24);
   B_25 : GTECH_BUF port map( A => N673, Z => N25);
   I_58 : GTECH_NOT port map( A => N263, Z => N264);
   C1943_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 3 )
      port map(
         -- Connections to port 'DATA1'
         DATA(2) => X_Logic0_port, DATA(1) => X_Logic1_port, DATA(0) => 
               X_Logic1_port, 
         -- Connections to port 'DATA2'
         DATA(5) => N262, DATA(4) => N261, DATA(3) => N260, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N18, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N19, 
         -- Connections to port 'Z'
         Z(2) => N267, Z(1) => N266, Z(0) => N265 );
   C1944_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => N661, 
         -- Connections to port 'DATA2'
         DATA(1) => X_Logic1_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N18, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N19, 
         -- Connections to port 'Z'
         Z(0) => N268 );
   C1945_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 2 )
      port map(
         -- Connections to port 'DATA1'
         DATA(1) => N259, DATA(0) => N258, 
         -- Connections to port 'DATA2'
         DATA(3) => N263, DATA(2) => N264, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N18, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N19, 
         -- Connections to port 'Z'
         Z(1) => N270, Z(0) => N269 );
   C1946_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 3 )
      port map(
         -- Connections to port 'DATA1'
         DATA(2) => X_Logic0_port, DATA(1) => X_Logic1_port, DATA(0) => 
               X_Logic1_port, 
         -- Connections to port 'DATA2'
         DATA(5) => cyc_s_2_port, DATA(4) => cyc_s_1_port, DATA(3) => 
               cyc_s_0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N20, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N230, 
         -- Connections to port 'Z'
         Z(2) => N273, Z(1) => N272, Z(0) => N271 );
   C1947_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 2 )
      port map(
         -- Connections to port 'DATA1'
         DATA(1) => N270, DATA(0) => N269, 
         -- Connections to port 'DATA2'
         DATA(3) => X_Logic0_port, DATA(2) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N26, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N253, 
         -- Connections to port 'Z'
         Z(1) => N275, Z(0) => N274 );
   B_26 : GTECH_BUF port map( A => N252, Z => N26);
   C1948_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 3 )
      port map(
         -- Connections to port 'DATA1'
         DATA(2) => N267, DATA(1) => N266, DATA(0) => N265, 
         -- Connections to port 'DATA2'
         DATA(5) => N273, DATA(4) => N272, DATA(3) => N271, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N26, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N253, 
         -- Connections to port 'Z'
         Z(2) => N278, Z(1) => N277, Z(0) => N276 );
   C1949_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => N268, 
         -- Connections to port 'DATA2'
         DATA(1) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N26, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N253, 
         -- Connections to port 'Z'
         Z(0) => N279 );
   C1950_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 2 )
      port map(
         -- Connections to port 'DATA1'
         DATA(1) => N275, DATA(0) => N274, 
         -- Connections to port 'DATA2'
         DATA(3) => X_Logic0_port, DATA(2) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N27, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N250, 
         -- Connections to port 'Z'
         Z(1) => N281, Z(0) => N280 );
   B_27 : GTECH_BUF port map( A => N249, Z => N27);
   C1951_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 3 )
      port map(
         -- Connections to port 'DATA1'
         DATA(2) => N278, DATA(1) => N277, DATA(0) => N276, 
         -- Connections to port 'DATA2'
         DATA(5) => X_Logic0_port, DATA(4) => X_Logic1_port, DATA(3) => 
               X_Logic1_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N27, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N250, 
         -- Connections to port 'Z'
         Z(2) => N284, Z(1) => N283, Z(0) => N282 );
   C1952_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => N279, 
         -- Connections to port 'DATA2'
         DATA(1) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N27, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N250, 
         -- Connections to port 'Z'
         Z(0) => N285 );
   C1953_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => N241, 
         -- Connections to port 'DATA2'
         DATA(1) => N285, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N28, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N187, 
         -- Connections to port 'Z'
         Z(0) => N286 );
   B_28 : GTECH_BUF port map( A => N186, Z => N28);
   C1954_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 2 )
      port map(
         -- Connections to port 'DATA1'
         DATA(1) => N243, DATA(0) => N242, 
         -- Connections to port 'DATA2'
         DATA(3) => N281, DATA(2) => N280, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N28, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N187, 
         -- Connections to port 'Z'
         Z(1) => N288, Z(0) => N287 );
   C1955_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 3 )
      port map(
         -- Connections to port 'DATA1'
         DATA(2) => N246, DATA(1) => N245, DATA(0) => N244, 
         -- Connections to port 'DATA2'
         DATA(5) => N284, DATA(4) => N283, DATA(3) => N282, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N28, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N187, 
         -- Connections to port 'Z'
         Z(2) => N291, Z(1) => N290, Z(0) => N289 );
   C1956_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => N247, 
         -- Connections to port 'DATA2'
         DATA(1) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N28, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N187, 
         -- Connections to port 'Z'
         Z(0) => N292 );
   C1957_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => N624, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N28, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N187, 
         -- Connections to port 'Z'
         Z(0) => N293 );
   C1958_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => N630, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N28, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N187, 
         -- Connections to port 'Z'
         Z(0) => N294 );
   C1959_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => N285, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N28, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N187, 
         -- Connections to port 'Z'
         Z(0) => N295 );
   C1960_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 3 )
      port map(
         -- Connections to port 'DATA1'
         DATA(2) => X_Logic0_port, DATA(1) => X_Logic1_port, DATA(0) => 
               X_Logic1_port, 
         -- Connections to port 'DATA2'
         DATA(5) => N291, DATA(4) => N290, DATA(3) => N289, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N29, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N184, 
         -- Connections to port 'Z'
         Z(2) => N298, Z(1) => N297, Z(0) => N296 );
   B_29 : GTECH_BUF port map( A => N183, Z => N29);
   C1961_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => N295, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N29, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N184, 
         -- Connections to port 'Z'
         Z(0) => N299 );
   C1962_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => N286, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N29, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N184, 
         -- Connections to port 'Z'
         Z(0) => N300 );
   C1963_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 2 )
      port map(
         -- Connections to port 'DATA1'
         DATA(1) => X_Logic0_port, DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(3) => N288, DATA(2) => N287, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N29, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N184, 
         -- Connections to port 'Z'
         Z(1) => N302, Z(0) => N301 );
   C1964_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => N292, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N29, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N184, 
         -- Connections to port 'Z'
         Z(0) => N303 );
   C1965_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => N293, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N29, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N184, 
         -- Connections to port 'Z'
         Z(0) => N304 );
   C1966_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => N294, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N29, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N184, 
         -- Connections to port 'Z'
         Z(0) => N305 );
   C1967_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => decrypt_in_port, 
         -- Connections to port 'DATA2'
         DATA(1) => decrypt_op_s, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N30, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N31, 
         -- Connections to port 'Z'
         Z(0) => N306 );
   B_30 : GTECH_BUF port map( A => N750, Z => N30);
   B_31 : GTECH_BUF port map( A => N749, Z => N31);
   C1968_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 3 )
      port map(
         -- Connections to port 'DATA1'
         DATA(2) => N181, DATA(1) => N180, DATA(0) => N179, 
         -- Connections to port 'DATA2'
         DATA(5) => N298, DATA(4) => N297, DATA(3) => N296, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N30, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N31, 
         -- Connections to port 'Z'
         Z(2) => N309, Z(1) => N308, Z(0) => N307 );
   C1969_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => bdi_valid_port, 
         -- Connections to port 'DATA2'
         DATA(1) => N300, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N30, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N31, 
         -- Connections to port 'Z'
         Z(0) => N310 );
   C1970_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 2 )
      port map(
         -- Connections to port 'DATA1'
         DATA(1) => X_Logic0_port, DATA(0) => bdi_valid_port, 
         -- Connections to port 'DATA2'
         DATA(3) => N302, DATA(2) => N301, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N30, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N31, 
         -- Connections to port 'Z'
         Z(1) => N312, Z(0) => N311 );
   C1971_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => N305, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N30, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N31, 
         -- Connections to port 'Z'
         Z(0) => N313 );
   C1972_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => N299, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N30, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N31, 
         -- Connections to port 'Z'
         Z(0) => N314 );
   C1973_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => N303, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N30, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N31, 
         -- Connections to port 'Z'
         Z(0) => N315 );
   C1974_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => N304, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N30, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N31, 
         -- Connections to port 'Z'
         Z(0) => N316 );
   I_59 : GTECH_NOT port map( A => N325, Z => N326);
   C1976_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 2 )
      port map(
         -- Connections to port 'DATA1'
         DATA(1) => X_Logic0_port, DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(3) => N325, DATA(2) => N326, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N32, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N324, 
         -- Connections to port 'Z'
         Z(1) => N328, Z(0) => N327 );
   B_32 : GTECH_BUF port map( A => N323, Z => N32);
   C1977_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 3 )
      port map(
         -- Connections to port 'DATA1'
         DATA(2) => X_Logic0_port, DATA(1) => X_Logic1_port, DATA(0) => 
               X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(5) => calling_state_2_port, DATA(4) => calling_state_1_port, 
               DATA(3) => calling_state_0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N18, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N19, 
         -- Connections to port 'Z'
         Z(2) => N334, Z(1) => N333, Z(0) => N332 );
   C1978_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => gtr_one_perm, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N18, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N19, 
         -- Connections to port 'Z'
         Z(0) => N335 );
   C1979_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => N753, 
         -- Connections to port 'DATA2'
         DATA(1) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N18, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N19, 
         -- Connections to port 'Z'
         Z(0) => N336 );
   C1980_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic1_port, 
         -- Connections to port 'DATA2'
         DATA(1) => gtr_one_perm, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N33, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N34, 
         -- Connections to port 'Z'
         Z(0) => N337 );
   B_33 : GTECH_BUF port map( A => N670, Z => N33);
   B_34 : GTECH_BUF port map( A => N669, Z => N34);
   C1981_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => N753, 
         -- Connections to port 'DATA2'
         DATA(1) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N33, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N34, 
         -- Connections to port 'Z'
         Z(0) => N338 );
   C1982_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 2 )
      port map(
         -- Connections to port 'DATA1'
         DATA(1) => bdi_size_1_port, DATA(0) => bdi_size_0_port, 
         -- Connections to port 'DATA2'
         DATA(3) => X_Logic0_port, DATA(2) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N35, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N331, 
         -- Connections to port 'Z'
         Z(1) => N340, Z(0) => N339 );
   B_35 : GTECH_BUF port map( A => N330, Z => N35);
   C1983_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 2 )
      port map(
         -- Connections to port 'DATA1'
         DATA(1) => bdi_eot_port, DATA(0) => N336, 
         -- Connections to port 'DATA2'
         DATA(3) => X_Logic0_port, DATA(2) => N338, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N35, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N331, 
         -- Connections to port 'Z'
         Z(1) => N342, Z(0) => N341 );
   C1984_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 3 )
      port map(
         -- Connections to port 'DATA1'
         DATA(2) => N334, DATA(1) => N333, DATA(0) => N332, 
         -- Connections to port 'DATA2'
         DATA(5) => calling_state_2_port, DATA(4) => calling_state_1_port, 
               DATA(3) => calling_state_0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N35, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N331, 
         -- Connections to port 'Z'
         Z(2) => N345, Z(1) => N344, Z(0) => N343 );
   C1985_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => N335, 
         -- Connections to port 'DATA2'
         DATA(1) => N337, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N35, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N331, 
         -- Connections to port 'Z'
         Z(0) => N346 );
   C1986_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 3 )
      port map(
         -- Connections to port 'DATA1'
         DATA(2) => X_Logic0_port, DATA(1) => X_Logic1_port, DATA(0) => 
               X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(5) => N345, DATA(4) => N344, DATA(3) => N343, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N36, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N37, 
         -- Connections to port 'Z'
         Z(2) => N349, Z(1) => N348, Z(0) => N347 );
   B_36 : GTECH_BUF port map( A => N721, Z => N36);
   B_37 : GTECH_BUF port map( A => N722, Z => N37);
   C1987_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => N346, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N36, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N37, 
         -- Connections to port 'Z'
         Z(0) => N350 );
   C1988_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 2 )
      port map(
         -- Connections to port 'DATA1'
         DATA(1) => X_Logic1_port, DATA(0) => N753, 
         -- Connections to port 'DATA2'
         DATA(3) => N342, DATA(2) => N341, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N36, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N37, 
         -- Connections to port 'Z'
         Z(1) => N352, Z(0) => N351 );
   C1989_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => N330, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N36, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N37, 
         -- Connections to port 'Z'
         Z(0) => N353 );
   C1990_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 2 )
      port map(
         -- Connections to port 'DATA1'
         DATA(1) => X_Logic0_port, DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(3) => N340, DATA(2) => N339, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N36, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N37, 
         -- Connections to port 'Z'
         Z(1) => N355, Z(0) => N354 );
   I_60 : GTECH_NOT port map( A => N360, Z => N361);
   C1992_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => N665, 
         -- Connections to port 'DATA2'
         DATA(1) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N0, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N1, 
         -- Connections to port 'Z'
         Z(0) => N367 );
   C1993_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => N624, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N0, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N1, 
         -- Connections to port 'Z'
         Z(0) => N368 );
   I_61 : GTECH_NOT port map( A => N369, Z => N370);
   I_62 : GTECH_NOT port map( A => N371, Z => N372);
   C1996_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => gtr_one_perm, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N18, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N19, 
         -- Connections to port 'Z'
         Z(0) => N373 );
   C1997_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 3 )
      port map(
         -- Connections to port 'DATA1'
         DATA(2) => X_Logic0_port, DATA(1) => X_Logic1_port, DATA(0) => 
               X_Logic1_port, 
         -- Connections to port 'DATA2'
         DATA(5) => calling_state_2_port, DATA(4) => calling_state_1_port, 
               DATA(3) => calling_state_0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N18, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N19, 
         -- Connections to port 'Z'
         Z(2) => N376, Z(1) => N375, Z(0) => N374 );
   C1998_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 2 )
      port map(
         -- Connections to port 'DATA1'
         DATA(1) => N369, DATA(0) => N370, 
         -- Connections to port 'DATA2'
         DATA(3) => N371, DATA(2) => N372, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N18, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N19, 
         -- Connections to port 'Z'
         Z(1) => N378, Z(0) => N377 );
   C1999_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 2 )
      port map(
         -- Connections to port 'DATA1'
         DATA(1) => bdi_size_1_port, DATA(0) => bdi_size_0_port, 
         -- Connections to port 'DATA2'
         DATA(3) => X_Logic0_port, DATA(2) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N38, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N365, 
         -- Connections to port 'Z'
         Z(1) => N380, Z(0) => N379 );
   B_38 : GTECH_BUF port map( A => N364, Z => N38);
   C2000_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => N368, 
         -- Connections to port 'DATA2'
         DATA(1) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N38, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N365, 
         -- Connections to port 'Z'
         Z(0) => N381 );
   C2001_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => N640, 
         -- Connections to port 'DATA2'
         DATA(1) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N38, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N365, 
         -- Connections to port 'Z'
         Z(0) => N382 );
   C2002_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => N367, 
         -- Connections to port 'DATA2'
         DATA(1) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N38, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N365, 
         -- Connections to port 'Z'
         Z(0) => N383 );
   C2003_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 3 )
      port map(
         -- Connections to port 'DATA1'
         DATA(2) => bdi_eot_port, DATA(1) => N378, DATA(0) => N377, 
         -- Connections to port 'DATA2'
         DATA(5) => X_Logic0_port, DATA(4) => N790, DATA(3) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N38, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N365, 
         -- Connections to port 'Z'
         Z(2) => N386, Z(1) => N385, Z(0) => N384 );
   C2004_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => N373, 
         -- Connections to port 'DATA2'
         DATA(1) => gtr_one_perm, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N38, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N365, 
         -- Connections to port 'Z'
         Z(0) => N387 );
   C2005_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 3 )
      port map(
         -- Connections to port 'DATA1'
         DATA(2) => N376, DATA(1) => N375, DATA(0) => N374, 
         -- Connections to port 'DATA2'
         DATA(5) => calling_state_2_port, DATA(4) => calling_state_1_port, 
               DATA(3) => calling_state_0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N38, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N365, 
         -- Connections to port 'Z'
         Z(2) => N390, Z(1) => N389, Z(0) => N388 );
   C2006_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 3 )
      port map(
         -- Connections to port 'DATA1'
         DATA(2) => X_Logic0_port, DATA(1) => X_Logic1_port, DATA(0) => 
               X_Logic1_port, 
         -- Connections to port 'DATA2'
         DATA(5) => N390, DATA(4) => N389, DATA(3) => N388, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N39, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N359, 
         -- Connections to port 'Z'
         Z(2) => N393, Z(1) => N392, Z(0) => N391 );
   B_39 : GTECH_BUF port map( A => N358, Z => N39);
   C2007_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => N387, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N39, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N359, 
         -- Connections to port 'Z'
         Z(0) => N394 );
   C2008_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 3 )
      port map(
         -- Connections to port 'DATA1'
         DATA(2) => X_Logic1_port, DATA(1) => N360, DATA(0) => N361, 
         -- Connections to port 'DATA2'
         DATA(5) => N386, DATA(4) => N385, DATA(3) => N384, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N39, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N359, 
         -- Connections to port 'Z'
         Z(2) => N397, Z(1) => N396, Z(0) => N395 );
   C2009_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => N364, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N39, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N359, 
         -- Connections to port 'Z'
         Z(0) => N398 );
   C2010_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 2 )
      port map(
         -- Connections to port 'DATA1'
         DATA(1) => X_Logic0_port, DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(3) => N380, DATA(2) => N379, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N39, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N359, 
         -- Connections to port 'Z'
         Z(1) => N400, Z(0) => N399 );
   C2011_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => N381, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N39, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N359, 
         -- Connections to port 'Z'
         Z(0) => N401 );
   C2012_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => N382, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N39, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N359, 
         -- Connections to port 'Z'
         Z(0) => N402 );
   C2013_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => N383, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N39, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N359, 
         -- Connections to port 'Z'
         Z(0) => N403 );
   I_63 : GTECH_NOT port map( A => N794, Z => N404);
   I_64 : GTECH_NOT port map( A => N798, Z => N405);
   C2016_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 2 )
      port map(
         -- Connections to port 'DATA1'
         DATA(1) => N404, DATA(0) => N794, 
         -- Connections to port 'DATA2'
         DATA(3) => N405, DATA(2) => N798, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N40, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N41, 
         -- Connections to port 'Z'
         Z(1) => N407, Z(0) => N406 );
   B_40 : GTECH_BUF port map( A => N753, Z => N40);
   B_41 : GTECH_BUF port map( A => gtr_one_perm, Z => N41);
   C2017_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 3 )
      port map(
         -- Connections to port 'DATA1'
         DATA(2) => X_Logic0_port, DATA(1) => X_Logic1_port, DATA(0) => 
               X_Logic1_port, 
         -- Connections to port 'DATA2'
         DATA(5) => calling_state_2_port, DATA(4) => calling_state_1_port, 
               DATA(3) => calling_state_0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N18, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N19, 
         -- Connections to port 'Z'
         Z(2) => N412, Z(1) => N411, Z(0) => N410 );
   C2018_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 2 )
      port map(
         -- Connections to port 'DATA1'
         DATA(1) => bdi_size_1_port, DATA(0) => bdi_size_0_port, 
         -- Connections to port 'DATA2'
         DATA(3) => X_Logic0_port, DATA(2) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N42, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N409, 
         -- Connections to port 'Z'
         Z(1) => N414, Z(0) => N413 );
   B_42 : GTECH_BUF port map( A => N408, Z => N42);
   C2019_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 3 )
      port map(
         -- Connections to port 'DATA1'
         DATA(2) => N412, DATA(1) => N411, DATA(0) => N410, 
         -- Connections to port 'DATA2'
         DATA(5) => calling_state_2_port, DATA(4) => calling_state_1_port, 
               DATA(3) => calling_state_0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N42, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N409, 
         -- Connections to port 'Z'
         Z(2) => N417, Z(1) => N416, Z(0) => N415 );
   C2020_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => gtr_one_perm, 
         -- Connections to port 'DATA2'
         DATA(1) => X_Logic1_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N42, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N409, 
         -- Connections to port 'Z'
         Z(0) => N418 );
   C2021_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => N418, 
         -- Connections to port 'DATA2'
         DATA(1) => gtr_one_perm, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N43, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N44, 
         -- Connections to port 'Z'
         Z(0) => N419 );
   B_43 : GTECH_BUF port map( A => N728, Z => N43);
   B_44 : GTECH_BUF port map( A => N727, Z => N44);
   C2022_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => N408, 
         -- Connections to port 'DATA2'
         DATA(1) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N43, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N44, 
         -- Connections to port 'Z'
         Z(0) => N420 );
   C2023_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 2 )
      port map(
         -- Connections to port 'DATA1'
         DATA(1) => N414, DATA(0) => N413, 
         -- Connections to port 'DATA2'
         DATA(3) => X_Logic0_port, DATA(2) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N43, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N44, 
         -- Connections to port 'Z'
         Z(1) => N422, Z(0) => N421 );
   C2024_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 3 )
      port map(
         -- Connections to port 'DATA1'
         DATA(2) => N417, DATA(1) => N416, DATA(0) => N415, 
         -- Connections to port 'DATA2'
         DATA(5) => X_Logic0_port, DATA(4) => X_Logic1_port, DATA(3) => 
               X_Logic1_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N43, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N44, 
         -- Connections to port 'Z'
         Z(2) => N425, Z(1) => N424, Z(0) => N423 );
   C2025_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 3 )
      port map(
         -- Connections to port 'DATA1'
         DATA(2) => N753, DATA(1) => N407, DATA(0) => N406, 
         -- Connections to port 'DATA2'
         DATA(5) => X_Logic0_port, DATA(4) => X_Logic0_port, DATA(3) => N801, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N45, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N46, 
         -- Connections to port 'Z'
         Z(2) => N428, Z(1) => N427, Z(0) => N426 );
   B_45 : GTECH_BUF port map( A => N718, Z => N45);
   B_46 : GTECH_BUF port map( A => N717, Z => N46);
   C2026_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => N753, 
         -- Connections to port 'DATA2'
         DATA(1) => N801, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N45, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N46, 
         -- Connections to port 'Z'
         Z(0) => N429 );
   C2027_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 3 )
      port map(
         -- Connections to port 'DATA1'
         DATA(2) => N425, DATA(1) => N424, DATA(0) => N423, 
         -- Connections to port 'DATA2'
         DATA(5) => calling_state_2_port, DATA(4) => calling_state_1_port, 
               DATA(3) => calling_state_0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N45, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N46, 
         -- Connections to port 'Z'
         Z(2) => N432, Z(1) => N431, Z(0) => N430 );
   C2028_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => N419, 
         -- Connections to port 'DATA2'
         DATA(1) => gtr_one_perm, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N45, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N46, 
         -- Connections to port 'Z'
         Z(0) => N433 );
   C2029_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => N420, 
         -- Connections to port 'DATA2'
         DATA(1) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N45, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N46, 
         -- Connections to port 'Z'
         Z(0) => N434 );
   C2030_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 2 )
      port map(
         -- Connections to port 'DATA1'
         DATA(1) => N422, DATA(0) => N421, 
         -- Connections to port 'DATA2'
         DATA(3) => X_Logic0_port, DATA(2) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N45, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N46, 
         -- Connections to port 'Z'
         Z(1) => N436, Z(0) => N435 );
   C2031_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => N403, 
         -- Connections to port 'DATA2'
         DATA(1) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N47, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N48, 
         -- Connections to port 'Z'
         Z(0) => N437 );
   B_47 : GTECH_BUF port map( A => N731, Z => N47);
   B_48 : GTECH_BUF port map( A => N730, Z => N48);
   C2032_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 3 )
      port map(
         -- Connections to port 'DATA1'
         DATA(2) => N393, DATA(1) => N392, DATA(0) => N391, 
         -- Connections to port 'DATA2'
         DATA(5) => N432, DATA(4) => N431, DATA(3) => N430, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N47, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N48, 
         -- Connections to port 'Z'
         Z(2) => N440, Z(1) => N439, Z(0) => N438 );
   C2033_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => N394, 
         -- Connections to port 'DATA2'
         DATA(1) => N433, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N47, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N48, 
         -- Connections to port 'Z'
         Z(0) => N441 );
   C2034_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 2 )
      port map(
         -- Connections to port 'DATA1'
         DATA(1) => N397, DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(3) => X_Logic0_port, DATA(2) => N429, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N47, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N48, 
         -- Connections to port 'Z'
         Z(1) => N443, Z(0) => N442 );
   C2035_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 3 )
      port map(
         -- Connections to port 'DATA1'
         DATA(2) => N397, DATA(1) => N396, DATA(0) => N395, 
         -- Connections to port 'DATA2'
         DATA(5) => N428, DATA(4) => N427, DATA(3) => N426, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N47, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N48, 
         -- Connections to port 'Z'
         Z(2) => N446, Z(1) => N445, Z(0) => N444 );
   C2036_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => N398, 
         -- Connections to port 'DATA2'
         DATA(1) => N434, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N47, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N48, 
         -- Connections to port 'Z'
         Z(0) => N447 );
   C2037_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 2 )
      port map(
         -- Connections to port 'DATA1'
         DATA(1) => N400, DATA(0) => N399, 
         -- Connections to port 'DATA2'
         DATA(3) => N436, DATA(2) => N435, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N47, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N48, 
         -- Connections to port 'Z'
         Z(1) => N449, Z(0) => N448 );
   C2038_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => N401, 
         -- Connections to port 'DATA2'
         DATA(1) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N47, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N48, 
         -- Connections to port 'Z'
         Z(0) => N450 );
   C2039_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => N402, 
         -- Connections to port 'DATA2'
         DATA(1) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N47, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N48, 
         -- Connections to port 'Z'
         Z(0) => N451 );
   C2040_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => N323, 
         -- Connections to port 'DATA2'
         DATA(1) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N49, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N50, 
         -- Connections to port 'Z'
         Z(0) => N452 );
   B_49 : GTECH_BUF port map( A => N740, Z => N49);
   B_50 : GTECH_BUF port map( A => N739, Z => N50);
   C2041_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 3 )
      port map(
         -- Connections to port 'DATA1'
         DATA(2) => X_Logic1_port, DATA(1) => N328, DATA(0) => N327, 
         -- Connections to port 'DATA2'
         DATA(5) => N446, DATA(4) => N445, DATA(3) => N444, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N49, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N50, 
         -- Connections to port 'Z'
         Z(2) => N455, Z(1) => N454, Z(0) => N453 );
   C2042_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 2 )
      port map(
         -- Connections to port 'DATA1'
         DATA(1) => N355, DATA(0) => N354, 
         -- Connections to port 'DATA2'
         DATA(3) => N449, DATA(2) => N448, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N49, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N50, 
         -- Connections to port 'Z'
         Z(1) => N457, Z(0) => N456 );
   C2043_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 3 )
      port map(
         -- Connections to port 'DATA1'
         DATA(2) => N349, DATA(1) => N348, DATA(0) => N347, 
         -- Connections to port 'DATA2'
         DATA(5) => N440, DATA(4) => N439, DATA(3) => N438, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N49, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N50, 
         -- Connections to port 'Z'
         Z(2) => N460, Z(1) => N459, Z(0) => N458 );
   C2044_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => N350, 
         -- Connections to port 'DATA2'
         DATA(1) => N441, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N49, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N50, 
         -- Connections to port 'Z'
         Z(0) => N461 );
   C2045_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 4 )
      port map(
         -- Connections to port 'DATA1'
         DATA(3) => N352, DATA(2) => X_Logic0_port, DATA(1) => N351, DATA(0) =>
               N351, 
         -- Connections to port 'DATA2'
         DATA(7) => X_Logic0_port, DATA(6) => N443, DATA(5) => X_Logic0_port, 
               DATA(4) => N442, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N49, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N50, 
         -- Connections to port 'Z'
         Z(3) => N465, Z(2) => N464, Z(1) => N463, Z(0) => N462 );
   C2046_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => N353, 
         -- Connections to port 'DATA2'
         DATA(1) => N447, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N49, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N50, 
         -- Connections to port 'Z'
         Z(0) => N466 );
   C2047_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => N451, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N49, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N50, 
         -- Connections to port 'Z'
         Z(0) => N467 );
   C2048_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => N437, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N49, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N50, 
         -- Connections to port 'Z'
         Z(0) => N468 );
   C2049_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => N450, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N49, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N50, 
         -- Connections to port 'Z'
         Z(0) => N469 );
   C2050_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 3 )
      port map(
         -- Connections to port 'DATA1'
         DATA(2) => X_Logic0_port, DATA(1) => X_Logic0_port, DATA(0) => 
               X_Logic1_port, 
         -- Connections to port 'DATA2'
         DATA(5) => N460, DATA(4) => N459, DATA(3) => N458, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N51, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N52, 
         -- Connections to port 'Z'
         Z(2) => N472, Z(1) => N471, Z(0) => N470 );
   B_51 : GTECH_BUF port map( A => N743, Z => N51);
   B_52 : GTECH_BUF port map( A => N742, Z => N52);
   C2051_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 4 )
      port map(
         -- Connections to port 'DATA1'
         DATA(3) => X_Logic0_port, DATA(2) => X_Logic0_port, DATA(1) => 
               X_Logic1_port, DATA(0) => X_Logic1_port, 
         -- Connections to port 'DATA2'
         DATA(7) => N465, DATA(6) => N464, DATA(5) => N463, DATA(4) => N462, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N51, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N52, 
         -- Connections to port 'Z'
         Z(3) => N476, Z(2) => N475, Z(1) => N474, Z(0) => N473 );
   C2052_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 3 )
      port map(
         -- Connections to port 'DATA1'
         DATA(2) => X_Logic1_port, DATA(1) => X_Logic1_port, DATA(0) => 
               X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(5) => N455, DATA(4) => N454, DATA(3) => N453, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N51, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N52, 
         -- Connections to port 'Z'
         Z(2) => N479, Z(1) => N478, Z(0) => N477 );
   C2053_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => N469, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N51, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N52, 
         -- Connections to port 'Z'
         Z(0) => N480 );
   C2054_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => N452, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N51, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N52, 
         -- Connections to port 'Z'
         Z(0) => N481 );
   C2055_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 2 )
      port map(
         -- Connections to port 'DATA1'
         DATA(1) => X_Logic0_port, DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(3) => N457, DATA(2) => N456, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N51, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N52, 
         -- Connections to port 'Z'
         Z(1) => N483, Z(0) => N482 );
   C2056_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => gtr_one_perm, 
         -- Connections to port 'DATA2'
         DATA(1) => N461, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N51, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N52, 
         -- Connections to port 'Z'
         Z(0) => N484 );
   C2057_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => N466, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N51, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N52, 
         -- Connections to port 'Z'
         Z(0) => N485 );
   C2058_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => N467, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N51, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N52, 
         -- Connections to port 'Z'
         Z(0) => N486 );
   C2059_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => N468, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N51, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N52, 
         -- Connections to port 'Z'
         Z(0) => N487 );
   I_65 : GTECH_NOT port map( A => N318, Z => N488);
   C2061_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 3 )
      port map(
         -- Connections to port 'DATA1'
         DATA(2) => cyc_s_2_port, DATA(1) => cyc_s_1_port, DATA(0) => 
               cyc_s_0_port, 
         -- Connections to port 'DATA2'
         DATA(5) => X_Logic1_port, DATA(4) => X_Logic0_port, DATA(3) => 
               X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N53, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N319, 
         -- Connections to port 'Z'
         Z(2) => N491, Z(1) => N490, Z(0) => N489 );
   B_53 : GTECH_BUF port map( A => N318, Z => N53);
   C2062_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => N487, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N53, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N319, 
         -- Connections to port 'Z'
         Z(0) => N492 );
   C2063_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 3 )
      port map(
         -- Connections to port 'DATA1'
         DATA(2) => calling_state_2_port, DATA(1) => calling_state_1_port, 
               DATA(0) => calling_state_0_port, 
         -- Connections to port 'DATA2'
         DATA(5) => N472, DATA(4) => N471, DATA(3) => N470, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N53, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N319, 
         -- Connections to port 'Z'
         Z(2) => N495, Z(1) => N494, Z(0) => N493 );
   C2064_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 4 )
      port map(
         -- Connections to port 'DATA1'
         DATA(3) => X_Logic0_port, DATA(2) => X_Logic0_port, DATA(1) => 
               X_Logic0_port, DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(7) => N476, DATA(6) => N475, DATA(5) => N474, DATA(4) => N473, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N53, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N319, 
         -- Connections to port 'Z'
         Z(3) => N499, Z(2) => N498, Z(1) => N497, Z(0) => N496 );
   C2065_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 3 )
      port map(
         -- Connections to port 'DATA1'
         DATA(2) => X_Logic0_port, DATA(1) => X_Logic0_port, DATA(0) => 
               X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(5) => N479, DATA(4) => N478, DATA(3) => N477, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N53, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N319, 
         -- Connections to port 'Z'
         Z(2) => N502, Z(1) => N501, Z(0) => N500 );
   C2066_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => N480, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N53, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N319, 
         -- Connections to port 'Z'
         Z(0) => N503 );
   C2067_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => N481, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N53, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N319, 
         -- Connections to port 'Z'
         Z(0) => N504 );
   C2068_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 2 )
      port map(
         -- Connections to port 'DATA1'
         DATA(1) => X_Logic0_port, DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(3) => N483, DATA(2) => N482, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N53, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N319, 
         -- Connections to port 'Z'
         Z(1) => N506, Z(0) => N505 );
   C2069_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => gtr_one_perm, 
         -- Connections to port 'DATA2'
         DATA(1) => N484, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N53, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N319, 
         -- Connections to port 'Z'
         Z(0) => N507 );
   C2070_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => N485, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N53, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N319, 
         -- Connections to port 'Z'
         Z(0) => N508 );
   C2071_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => N486, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N53, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N319, 
         -- Connections to port 'Z'
         Z(0) => N509 );
   C2072_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 3 )
      port map(
         -- Connections to port 'DATA1'
         DATA(2) => X_Logic0_port, DATA(1) => X_Logic0_port, DATA(0) => 
               X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(5) => calling_state_2_port, DATA(4) => calling_state_1_port, 
               DATA(3) => calling_state_0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N54, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N55, 
         -- Connections to port 'Z'
         Z(2) => N514, Z(1) => N513, Z(0) => N512 );
   B_54 : GTECH_BUF port map( A => N649, Z => N54);
   B_55 : GTECH_BUF port map( A => N648, Z => N55);
   I_66 : GTECH_NOT port map( A => N510, Z => N515);
   C2074_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => N649, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N56, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N511, 
         -- Connections to port 'Z'
         Z(0) => N516 );
   B_56 : GTECH_BUF port map( A => N510, Z => N56);
   C2075_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 3 )
      port map(
         -- Connections to port 'DATA1'
         DATA(2) => calling_state_2_port, DATA(1) => calling_state_1_port, 
               DATA(0) => calling_state_0_port, 
         -- Connections to port 'DATA2'
         DATA(5) => N514, DATA(4) => N513, DATA(3) => N512, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N56, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N511, 
         -- Connections to port 'Z'
         Z(2) => N519, Z(1) => N518, Z(0) => N517 );
   C2076_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 3 )
      port map(
         -- Connections to port 'DATA1'
         DATA(2) => N519, DATA(1) => N518, DATA(0) => N517, 
         -- Connections to port 'DATA2'
         DATA(5) => calling_state_2_port, DATA(4) => calling_state_1_port, 
               DATA(3) => calling_state_0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N57, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N58, 
         -- Connections to port 'Z'
         Z(2) => N522, Z(1) => N521, Z(0) => N520 );
   B_57 : GTECH_BUF port map( A => N706, Z => N57);
   B_58 : GTECH_BUF port map( A => N705, Z => N58);
   C2077_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 3 )
      port map(
         -- Connections to port 'DATA1'
         DATA(2) => N510, DATA(1) => N515, DATA(0) => N510, 
         -- Connections to port 'DATA2'
         DATA(5) => cyc_s_2_port, DATA(4) => cyc_s_1_port, DATA(3) => 
               cyc_s_0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N57, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N58, 
         -- Connections to port 'Z'
         Z(2) => N525, Z(1) => N524, Z(0) => N523 );
   C2078_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => N516, 
         -- Connections to port 'DATA2'
         DATA(1) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N57, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N58, 
         -- Connections to port 'Z'
         Z(0) => N526 );
   C2079_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 3 )
      port map(
         -- Connections to port 'DATA1'
         DATA(2) => X_Logic1_port, DATA(1) => X_Logic0_port, DATA(0) => 
               X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(5) => calling_state_2_port, DATA(4) => calling_state_1_port, 
               DATA(3) => calling_state_0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N59, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N529, 
         -- Connections to port 'Z'
         Z(2) => N532, Z(1) => N531, Z(0) => N530 );
   B_59 : GTECH_BUF port map( A => N528, Z => N59);
   I_67 : GTECH_NOT port map( A => N528, Z => N533);
   C2081_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => N533, 
         -- Connections to port 'DATA2'
         DATA(1) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N60, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N61, 
         -- Connections to port 'Z'
         Z(0) => N534 );
   B_60 : GTECH_BUF port map( A => N678, Z => N60);
   B_61 : GTECH_BUF port map( A => N677, Z => N61);
   C2082_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 3 )
      port map(
         -- Connections to port 'DATA1'
         DATA(2) => X_Logic0_port, DATA(1) => N528, DATA(0) => N528, 
         -- Connections to port 'DATA2'
         DATA(5) => cyc_s_2_port, DATA(4) => cyc_s_1_port, DATA(3) => 
               cyc_s_0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N60, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N61, 
         -- Connections to port 'Z'
         Z(2) => N537, Z(1) => N536, Z(0) => N535 );
   C2083_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 3 )
      port map(
         -- Connections to port 'DATA1'
         DATA(2) => N532, DATA(1) => N531, DATA(0) => N530, 
         -- Connections to port 'DATA2'
         DATA(5) => calling_state_2_port, DATA(4) => calling_state_1_port, 
               DATA(3) => calling_state_0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N60, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N61, 
         -- Connections to port 'Z'
         Z(2) => N540, Z(1) => N539, Z(0) => N538 );
   C2084_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => N528, 
         -- Connections to port 'DATA2'
         DATA(1) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N60, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N61, 
         -- Connections to port 'Z'
         Z(0) => N541 );
   C2085_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => tag_verified, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N62, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N547, 
         -- Connections to port 'Z'
         Z(0) => N548 );
   B_62 : GTECH_BUF port map( A => N546, Z => N62);
   I_68 : GTECH_NOT port map( A => N549, Z => N550);
   C2087_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 3 )
      port map(
         -- Connections to port 'DATA1'
         DATA(2) => X_Logic0_port, DATA(1) => X_Logic0_port, DATA(0) => 
               X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(5) => cyc_s_2_port, DATA(4) => cyc_s_1_port, DATA(3) => 
               cyc_s_0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N63, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N64, 
         -- Connections to port 'Z'
         Z(2) => N553, Z(1) => N552, Z(0) => N551 );
   B_63 : GTECH_BUF port map( A => N682, Z => N63);
   B_64 : GTECH_BUF port map( A => N681, Z => N64);
   C2088_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => N548, 
         -- Connections to port 'DATA2'
         DATA(1) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N63, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N64, 
         -- Connections to port 'Z'
         Z(0) => N554 );
   C2089_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic1_port, 
         -- Connections to port 'DATA2'
         DATA(1) => N550, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N63, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N64, 
         -- Connections to port 'Z'
         Z(0) => N555 );
   C2090_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => N555, 
         -- Connections to port 'DATA2'
         DATA(1) => X_Logic1_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N65, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N544, 
         -- Connections to port 'Z'
         Z(0) => N556 );
   B_65 : GTECH_BUF port map( A => N543, Z => N65);
   C2091_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => N682, 
         -- Connections to port 'DATA2'
         DATA(1) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N65, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N544, 
         -- Connections to port 'Z'
         Z(0) => N557 );
   C2092_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => N554, 
         -- Connections to port 'DATA2'
         DATA(1) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N65, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N544, 
         -- Connections to port 'Z'
         Z(0) => N558 );
   C2093_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 4 )
      port map(
         -- Connections to port 'DATA1'
         DATA(3) => X_Logic1_port, DATA(2) => X_Logic1_port, DATA(1) => 
               X_Logic1_port, DATA(0) => X_Logic1_port, 
         -- Connections to port 'DATA2'
         DATA(7) => bdi_valid_bytes_3_port, DATA(6) => bdi_valid_bytes_2_port, 
               DATA(5) => bdi_valid_bytes_1_port, DATA(4) => 
               bdi_valid_bytes_0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N66, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N67, 
         -- Connections to port 'Z'
         Z(3) => N562, Z(2) => N561, Z(1) => N560, Z(0) => N559 );
   B_66 : GTECH_BUF port map( A => N708, Z => N66);
   B_67 : GTECH_BUF port map( A => decrypt_op_s, Z => N67);
   C2094_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => bdo_ready_port, 
         -- Connections to port 'DATA2'
         DATA(1) => N543, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N66, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N67, 
         -- Connections to port 'Z'
         Z(0) => N563 );
   C2095_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => N541, 
         -- Connections to port 'DATA2'
         DATA(1) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N66, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N67, 
         -- Connections to port 'Z'
         Z(0) => N564 );
   C2096_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => N534, 
         -- Connections to port 'DATA2'
         DATA(1) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N66, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N67, 
         -- Connections to port 'Z'
         Z(0) => N565 );
   C2097_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 3 )
      port map(
         -- Connections to port 'DATA1'
         DATA(2) => N537, DATA(1) => N536, DATA(0) => N535, 
         -- Connections to port 'DATA2'
         DATA(5) => N553, DATA(4) => N552, DATA(3) => N551, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N66, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N67, 
         -- Connections to port 'Z'
         Z(2) => N568, Z(1) => N567, Z(0) => N566 );
   C2098_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => N558, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N66, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N67, 
         -- Connections to port 'Z'
         Z(0) => N569 );
   C2099_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => N543, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N66, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N67, 
         -- Connections to port 'Z'
         Z(0) => N570 );
   C2100_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic1_port, 
         -- Connections to port 'DATA2'
         DATA(1) => N556, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N66, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N67, 
         -- Connections to port 'Z'
         Z(0) => N571 );
   C2101_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => N557, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N66, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N67, 
         -- Connections to port 'Z'
         Z(0) => N572 );
   C2102_cell : SELECT_OP
      generic map ( num_inputs => 6, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => X_Logic1_port, 
         -- Connections to port 'DATA3'
         DATA(2) => X_Logic1_port, 
         -- Connections to port 'DATA4'
         DATA(3) => X_Logic1_port, 
         -- Connections to port 'DATA5'
         DATA(4) => X_Logic1_port, 
         -- Connections to port 'DATA6'
         DATA(5) => N571, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N68, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N69, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N70, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N71, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N72, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N73, 
         -- Connections to port 'Z'
         Z(0) => n_tag_verified );
   B_68 : GTECH_BUF port map( A => state_main_sel_5_port, Z => N68);
   B_69 : GTECH_BUF port map( A => N81, Z => N69);
   B_70 : GTECH_BUF port map( A => N84, Z => N70);
   B_71 : GTECH_BUF port map( A => N87, Z => N71);
   B_72 : GTECH_BUF port map( A => N90, Z => N72);
   B_73 : GTECH_BUF port map( A => N93, Z => N73);
   C2103_cell : SELECT_OP
      generic map ( num_inputs => 6, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic1_port, 
         -- Connections to port 'DATA2'
         DATA(1) => N173, 
         -- Connections to port 'DATA3'
         DATA(2) => X_Logic0_port, 
         -- Connections to port 'DATA4'
         DATA(3) => N488, 
         -- Connections to port 'DATA5'
         DATA(4) => N706, 
         -- Connections to port 'DATA6'
         DATA(5) => N564, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N68, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N69, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N70, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N71, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N72, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N73, 
         -- Connections to port 'Z'
         Z(0) => load_dcount );
   C2104_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => N507, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N68, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N71, 
         -- Connections to port 'Z'
         Z(0) => n_gtr_one_perm );
   C2105_cell : SELECT_OP
      generic map ( num_inputs => 6, input_width => 4 )
      port map(
         -- Connections to port 'DATA1'
         DATA(3) => X_Logic0_port, DATA(2) => N101, DATA(1) => N101, DATA(0) =>
               N101, 
         -- Connections to port 'DATA2'
         DATA(7) => X_Logic0_port, DATA(6) => X_Logic0_port, DATA(5) => 
               X_Logic0_port, DATA(4) => X_Logic0_port, 
         -- Connections to port 'DATA3'
         DATA(11) => N315, DATA(10) => X_Logic0_port, DATA(9) => X_Logic0_port,
               DATA(8) => X_Logic0_port, 
         -- Connections to port 'DATA4'
         DATA(15) => N504, DATA(14) => X_Logic0_port, DATA(13) => X_Logic0_port
               , DATA(12) => X_Logic0_port, 
         -- Connections to port 'DATA5'
         DATA(19) => X_Logic0_port, DATA(18) => X_Logic1_port, DATA(17) => 
               X_Logic1_port, DATA(16) => X_Logic1_port, 
         -- Connections to port 'DATA6'
         DATA(23) => X_Logic0_port, DATA(22) => X_Logic0_port, DATA(21) => 
               X_Logic0_port, DATA(20) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N68, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N69, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N70, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N71, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N72, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N73, 
         -- Connections to port 'Z'
         Z(3) => state_main_sel_6_port, Z(2) => state_main_sel_4_port, Z(1) => 
               state_main_sel_2, Z(0) => state_main_sel_0 );
   C2106_cell : SELECT_OP
      generic map ( num_inputs => 6, input_width => 3 )
      port map(
         -- Connections to port 'DATA1'
         DATA(2) => X_Logic1_port, DATA(1) => X_Logic1_port, DATA(0) => 
               X_Logic1_port, 
         -- Connections to port 'DATA2'
         DATA(5) => N173, DATA(4) => N173, DATA(3) => key_valid_port, 
         -- Connections to port 'DATA3'
         DATA(8) => N315, DATA(7) => N312, DATA(6) => N311, 
         -- Connections to port 'DATA4'
         DATA(11) => N502, DATA(10) => N501, DATA(9) => N500, 
         -- Connections to port 'DATA5'
         DATA(14) => X_Logic1_port, DATA(13) => X_Logic1_port, DATA(12) => 
               X_Logic1_port, 
         -- Connections to port 'DATA6'
         DATA(17) => X_Logic0_port, DATA(16) => X_Logic0_port, DATA(15) => 
               X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N68, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N69, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N70, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N71, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N72, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N73, 
         -- Connections to port 'Z'
         Z(2) => state_main_en_2_port, Z(1) => state_main_en_1_port, Z(0) => 
               state_main_en_0_port );
   C2107_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => N306, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N68, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N70, 
         -- Connections to port 'Z'
         Z(0) => n_decrypt_op_s );
   C2108_cell : SELECT_OP
      generic map ( num_inputs => 6, input_width => 3 )
      port map(
         -- Connections to port 'DATA1'
         DATA(2) => X_Logic0_port, DATA(1) => N99, DATA(0) => N98, 
         -- Connections to port 'DATA2'
         DATA(5) => N137, DATA(4) => N136, DATA(3) => N135, 
         -- Connections to port 'DATA3'
         DATA(8) => N309, DATA(7) => N308, DATA(6) => N307, 
         -- Connections to port 'DATA4'
         DATA(11) => N491, DATA(10) => N490, DATA(9) => N489, 
         -- Connections to port 'DATA5'
         DATA(14) => N525, DATA(13) => N524, DATA(12) => N523, 
         -- Connections to port 'DATA6'
         DATA(17) => N568, DATA(16) => N567, DATA(15) => N566, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N68, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N69, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N70, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N71, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N72, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N73, 
         -- Connections to port 'Z'
         Z(2) => n_cyc_s_2_port, Z(1) => n_cyc_s_1_port, Z(0) => n_cyc_s_0_port
               );
   C2109_cell : SELECT_OP
      generic map ( num_inputs => 5, input_width => 3 )
      port map(
         -- Connections to port 'DATA1'
         DATA(2) => hash_in_port, DATA(1) => X_Logic0_port, DATA(0) => 
               hash_in_port, 
         -- Connections to port 'DATA2'
         DATA(5) => N140, DATA(4) => N139, DATA(3) => N138, 
         -- Connections to port 'DATA3'
         DATA(8) => N495, DATA(7) => N494, DATA(6) => N493, 
         -- Connections to port 'DATA4'
         DATA(11) => N522, DATA(10) => N521, DATA(9) => N520, 
         -- Connections to port 'DATA5'
         DATA(14) => N540, DATA(13) => N539, DATA(12) => N538, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N68, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N69, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N71, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N72, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N73, 
         -- Connections to port 'Z'
         Z(2) => n_calling_state_2_port, Z(1) => n_calling_state_1_port, Z(0) 
               => n_calling_state_0_port );
   C2110_cell : SELECT_OP
      generic map ( num_inputs => 6, input_width => 32 )
      port map(
         -- Connections to port 'DATA1'
         DATA(31) => bdi_31_port, DATA(30) => bdi_30_port, DATA(29) => 
               bdi_29_port, DATA(28) => bdi_28_port, DATA(27) => bdi_27_port, 
               DATA(26) => bdi_26_port, DATA(25) => bdi_25_port, DATA(24) => 
               bdi_24_port, DATA(23) => bdi_23_port, DATA(22) => bdi_22_port, 
               DATA(21) => bdi_21_port, DATA(20) => bdi_20_port, DATA(19) => 
               bdi_19_port, DATA(18) => bdi_18_port, DATA(17) => bdi_17_port, 
               DATA(16) => bdi_16_port, DATA(15) => bdi_15_port, DATA(14) => 
               bdi_14_port, DATA(13) => bdi_13_port, DATA(12) => bdi_12_port, 
               DATA(11) => bdi_11_port, DATA(10) => bdi_10_port, DATA(9) => 
               bdi_9_port, DATA(8) => bdi_8_port, DATA(7) => bdi_7_port, 
               DATA(6) => bdi_6_port, DATA(5) => bdi_5_port, DATA(4) => 
               bdi_4_port, DATA(3) => bdi_3_port, DATA(2) => bdi_2_port, 
               DATA(1) => bdi_1_port, DATA(0) => bdi_0_port, 
         -- Connections to port 'DATA2'
         DATA(63) => N172, DATA(62) => N171, DATA(61) => N170, DATA(60) => N169
               , DATA(59) => N168, DATA(58) => N167, DATA(57) => N166, DATA(56)
               => N165, DATA(55) => N164, DATA(54) => N163, DATA(53) => N162, 
               DATA(52) => N161, DATA(51) => N160, DATA(50) => N159, DATA(49) 
               => N158, DATA(48) => N157, DATA(47) => N156, DATA(46) => N155, 
               DATA(45) => N154, DATA(44) => N153, DATA(43) => N152, DATA(42) 
               => N151, DATA(41) => N150, DATA(40) => N149, DATA(39) => N148, 
               DATA(38) => N147, DATA(37) => N146, DATA(36) => N145, DATA(35) 
               => N144, DATA(34) => N143, DATA(33) => N142, DATA(32) => N141, 
         -- Connections to port 'DATA3'
         DATA(95) => bdi_31_port, DATA(94) => bdi_30_port, DATA(93) => 
               bdi_29_port, DATA(92) => bdi_28_port, DATA(91) => bdi_27_port, 
               DATA(90) => bdi_26_port, DATA(89) => bdi_25_port, DATA(88) => 
               bdi_24_port, DATA(87) => bdi_23_port, DATA(86) => bdi_22_port, 
               DATA(85) => bdi_21_port, DATA(84) => bdi_20_port, DATA(83) => 
               bdi_19_port, DATA(82) => bdi_18_port, DATA(81) => bdi_17_port, 
               DATA(80) => bdi_16_port, DATA(79) => bdi_15_port, DATA(78) => 
               bdi_14_port, DATA(77) => bdi_13_port, DATA(76) => bdi_12_port, 
               DATA(75) => bdi_11_port, DATA(74) => bdi_10_port, DATA(73) => 
               bdi_9_port, DATA(72) => bdi_8_port, DATA(71) => bdi_7_port, 
               DATA(70) => bdi_6_port, DATA(69) => bdi_5_port, DATA(68) => 
               bdi_4_port, DATA(67) => bdi_3_port, DATA(66) => bdi_2_port, 
               DATA(65) => bdi_1_port, DATA(64) => bdi_0_port, 
         -- Connections to port 'DATA4'
         DATA(127) => bdi_31_port, DATA(126) => bdi_30_port, DATA(125) => 
               bdi_29_port, DATA(124) => bdi_28_port, DATA(123) => bdi_27_port,
               DATA(122) => bdi_26_port, DATA(121) => bdi_25_port, DATA(120) =>
               bdi_24_port, DATA(119) => bdi_23_port, DATA(118) => bdi_22_port,
               DATA(117) => bdi_21_port, DATA(116) => bdi_20_port, DATA(115) =>
               bdi_19_port, DATA(114) => bdi_18_port, DATA(113) => bdi_17_port,
               DATA(112) => bdi_16_port, DATA(111) => bdi_15_port, DATA(110) =>
               bdi_14_port, DATA(109) => bdi_13_port, DATA(108) => bdi_12_port,
               DATA(107) => bdi_11_port, DATA(106) => bdi_10_port, DATA(105) =>
               bdi_9_port, DATA(104) => bdi_8_port, DATA(103) => bdi_7_port, 
               DATA(102) => bdi_6_port, DATA(101) => bdi_5_port, DATA(100) => 
               bdi_4_port, DATA(99) => bdi_3_port, DATA(98) => bdi_2_port, 
               DATA(97) => bdi_1_port, DATA(96) => bdi_0_port, 
         -- Connections to port 'DATA5'
         DATA(159) => bdi_31_port, DATA(158) => bdi_30_port, DATA(157) => 
               bdi_29_port, DATA(156) => bdi_28_port, DATA(155) => bdi_27_port,
               DATA(154) => bdi_26_port, DATA(153) => bdi_25_port, DATA(152) =>
               bdi_24_port, DATA(151) => bdi_23_port, DATA(150) => bdi_22_port,
               DATA(149) => bdi_21_port, DATA(148) => bdi_20_port, DATA(147) =>
               bdi_19_port, DATA(146) => bdi_18_port, DATA(145) => bdi_17_port,
               DATA(144) => bdi_16_port, DATA(143) => bdi_15_port, DATA(142) =>
               bdi_14_port, DATA(141) => bdi_13_port, DATA(140) => bdi_12_port,
               DATA(139) => bdi_11_port, DATA(138) => bdi_10_port, DATA(137) =>
               bdi_9_port, DATA(136) => bdi_8_port, DATA(135) => bdi_7_port, 
               DATA(134) => bdi_6_port, DATA(133) => bdi_5_port, DATA(132) => 
               bdi_4_port, DATA(131) => bdi_3_port, DATA(130) => bdi_2_port, 
               DATA(129) => bdi_1_port, DATA(128) => bdi_0_port, 
         -- Connections to port 'DATA6'
         DATA(191) => bdi_31_port, DATA(190) => bdi_30_port, DATA(189) => 
               bdi_29_port, DATA(188) => bdi_28_port, DATA(187) => bdi_27_port,
               DATA(186) => bdi_26_port, DATA(185) => bdi_25_port, DATA(184) =>
               bdi_24_port, DATA(183) => bdi_23_port, DATA(182) => bdi_22_port,
               DATA(181) => bdi_21_port, DATA(180) => bdi_20_port, DATA(179) =>
               bdi_19_port, DATA(178) => bdi_18_port, DATA(177) => bdi_17_port,
               DATA(176) => bdi_16_port, DATA(175) => bdi_15_port, DATA(174) =>
               bdi_14_port, DATA(173) => bdi_13_port, DATA(172) => bdi_12_port,
               DATA(171) => bdi_11_port, DATA(170) => bdi_10_port, DATA(169) =>
               bdi_9_port, DATA(168) => bdi_8_port, DATA(167) => bdi_7_port, 
               DATA(166) => bdi_6_port, DATA(165) => bdi_5_port, DATA(164) => 
               bdi_4_port, DATA(163) => bdi_3_port, DATA(162) => bdi_2_port, 
               DATA(161) => bdi_1_port, DATA(160) => bdi_0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N68, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N69, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N70, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N71, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N72, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N73, 
         -- Connections to port 'Z'
         Z(31) => bdi_key_31_port, Z(30) => bdi_key_30_port, Z(29) => 
               bdi_key_29_port, Z(28) => bdi_key_28_port, Z(27) => 
               bdi_key_27_port, Z(26) => bdi_key_26_port, Z(25) => 
               bdi_key_25_port, Z(24) => bdi_key_24_port, Z(23) => 
               bdi_key_23_port, Z(22) => bdi_key_22_port, Z(21) => 
               bdi_key_21_port, Z(20) => bdi_key_20_port, Z(19) => 
               bdi_key_19_port, Z(18) => bdi_key_18_port, Z(17) => 
               bdi_key_17_port, Z(16) => bdi_key_16_port, Z(15) => 
               bdi_key_15_port, Z(14) => bdi_key_14_port, Z(13) => 
               bdi_key_13_port, Z(12) => bdi_key_12_port, Z(11) => 
               bdi_key_11_port, Z(10) => bdi_key_10_port, Z(9) => 
               bdi_key_9_port, Z(8) => bdi_key_8_port, Z(7) => bdi_key_7_port, 
               Z(6) => bdi_key_6_port, Z(5) => bdi_key_5_port, Z(4) => 
               bdi_key_4_port, Z(3) => bdi_key_3_port, Z(2) => bdi_key_2_port, 
               Z(1) => bdi_key_1_port, Z(0) => bdi_key_0_port );
   C2111_cell : SELECT_OP
      generic map ( num_inputs => 6, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => key_valid_port, 
         -- Connections to port 'DATA3'
         DATA(2) => X_Logic0_port, 
         -- Connections to port 'DATA4'
         DATA(3) => X_Logic0_port, 
         -- Connections to port 'DATA5'
         DATA(4) => X_Logic0_port, 
         -- Connections to port 'DATA6'
         DATA(5) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N68, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N69, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N70, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N71, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N72, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N73, 
         -- Connections to port 'Z'
         Z(0) => key_ready_port );
   C2112_cell : SELECT_OP
      generic map ( num_inputs => 6, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => key_valid_port, 
         -- Connections to port 'DATA3'
         DATA(2) => N310, 
         -- Connections to port 'DATA4'
         DATA(3) => N488, 
         -- Connections to port 'DATA5'
         DATA(4) => X_Logic0_port, 
         -- Connections to port 'DATA6'
         DATA(5) => N563, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N68, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N69, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N70, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N71, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N72, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N73, 
         -- Connections to port 'Z'
         Z(0) => en_dcount );
   C2113_cell : SELECT_OP
      generic map ( num_inputs => 6, input_width => 4 )
      port map(
         -- Connections to port 'DATA1'
         DATA(3) => X_Logic0_port, DATA(2) => X_Logic0_port, DATA(1) => 
               X_Logic0_port, DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(7) => X_Logic0_port, DATA(6) => X_Logic0_port, DATA(5) => N173, 
               DATA(4) => X_Logic0_port, 
         -- Connections to port 'DATA3'
         DATA(11) => X_Logic0_port, DATA(10) => X_Logic0_port, DATA(9) => 
               X_Logic0_port, DATA(8) => X_Logic0_port, 
         -- Connections to port 'DATA4'
         DATA(15) => N499, DATA(14) => N498, DATA(13) => N497, DATA(12) => N496
               , 
         -- Connections to port 'DATA5'
         DATA(19) => X_Logic0_port, DATA(18) => X_Logic0_port, DATA(17) => 
               X_Logic0_port, DATA(16) => X_Logic0_port, 
         -- Connections to port 'DATA6'
         DATA(23) => X_Logic0_port, DATA(22) => X_Logic0_port, DATA(21) => 
               X_Logic0_port, DATA(20) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N68, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N69, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N70, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N71, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N72, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N73, 
         -- Connections to port 'Z'
         Z(3) => cu_cd_s_7_port, Z(2) => cu_cd_s_6_port, Z(1) => cu_cd_s_1, 
               Z(0) => cu_cd_s_0 );
   C2114_cell : SELECT_OP
      generic map ( num_inputs => 6, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => N173, 
         -- Connections to port 'DATA3'
         DATA(2) => X_Logic0_port, 
         -- Connections to port 'DATA4'
         DATA(3) => N488, 
         -- Connections to port 'DATA5'
         DATA(4) => N706, 
         -- Connections to port 'DATA6'
         DATA(5) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N68, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N69, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N70, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N71, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N72, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N73, 
         -- Connections to port 'Z'
         Z(0) => load_rnd );
   C2115_cell : SELECT_OP
      generic map ( num_inputs => 6, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => X_Logic0_port, 
         -- Connections to port 'DATA3'
         DATA(2) => bdi_eot_port, 
         -- Connections to port 'DATA4'
         DATA(3) => X_Logic0_port, 
         -- Connections to port 'DATA5'
         DATA(4) => X_Logic0_port, 
         -- Connections to port 'DATA6'
         DATA(5) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N68, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N69, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N70, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N71, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N72, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N73, 
         -- Connections to port 'Z'
         Z(0) => n_bdi_eot_prev );
   C2116_cell : SELECT_OP
      generic map ( num_inputs => 6, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => X_Logic0_port, 
         -- Connections to port 'DATA3'
         DATA(2) => N316, 
         -- Connections to port 'DATA4'
         DATA(3) => N503, 
         -- Connections to port 'DATA5'
         DATA(4) => X_Logic0_port, 
         -- Connections to port 'DATA6'
         DATA(5) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N68, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N69, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N70, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N71, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N72, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N73, 
         -- Connections to port 'Z'
         Z(0) => cyc_state_update_sel );
   C2117_cell : SELECT_OP
      generic map ( num_inputs => 6, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => X_Logic0_port, 
         -- Connections to port 'DATA3'
         DATA(2) => N310, 
         -- Connections to port 'DATA4'
         DATA(3) => N508, 
         -- Connections to port 'DATA5'
         DATA(4) => X_Logic0_port, 
         -- Connections to port 'DATA6'
         DATA(5) => N570, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N68, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N69, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N70, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N71, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N72, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N73, 
         -- Connections to port 'Z'
         Z(0) => bdi_ready_port );
   C2118_cell : SELECT_OP
      generic map ( num_inputs => 6, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => X_Logic0_port, 
         -- Connections to port 'DATA3'
         DATA(2) => N313, 
         -- Connections to port 'DATA4'
         DATA(3) => N492, 
         -- Connections to port 'DATA5'
         DATA(4) => X_Logic0_port, 
         -- Connections to port 'DATA6'
         DATA(5) => N565, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N68, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N69, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N70, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N71, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N72, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N73, 
         -- Connections to port 'Z'
         Z(0) => end_of_block_port );
   C2119_cell : SELECT_OP
      generic map ( num_inputs => 6, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => X_Logic0_port, 
         -- Connections to port 'DATA3'
         DATA(2) => N314, 
         -- Connections to port 'DATA4'
         DATA(3) => N509, 
         -- Connections to port 'DATA5'
         DATA(4) => X_Logic0_port, 
         -- Connections to port 'DATA6'
         DATA(5) => N708, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N68, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N69, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N70, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N71, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N72, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N73, 
         -- Connections to port 'Z'
         Z(0) => bdo_valid_port );
   C2120_cell : SELECT_OP
      generic map ( num_inputs => 6, input_width => 2 )
      port map(
         -- Connections to port 'DATA1'
         DATA(1) => X_Logic0_port, DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(3) => X_Logic0_port, DATA(2) => X_Logic0_port, 
         -- Connections to port 'DATA3'
         DATA(5) => X_Logic0_port, DATA(4) => X_Logic0_port, 
         -- Connections to port 'DATA4'
         DATA(7) => N506, DATA(6) => N505, 
         -- Connections to port 'DATA5'
         DATA(9) => X_Logic0_port, DATA(8) => X_Logic0_port, 
         -- Connections to port 'DATA6'
         DATA(11) => X_Logic0_port, DATA(10) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N68, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N69, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N70, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N71, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N72, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N73, 
         -- Connections to port 'Z'
         Z(1) => cycd_sel_1_port, Z(0) => cycd_sel_0_port );
   C2121_cell : SELECT_OP
      generic map ( num_inputs => 6, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => X_Logic0_port, 
         -- Connections to port 'DATA3'
         DATA(2) => X_Logic0_port, 
         -- Connections to port 'DATA4'
         DATA(3) => X_Logic0_port, 
         -- Connections to port 'DATA5'
         DATA(4) => X_Logic1_port, 
         -- Connections to port 'DATA6'
         DATA(5) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N68, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N69, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N70, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N71, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N72, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N73, 
         -- Connections to port 'Z'
         Z(0) => en_rnd );
   C2122_cell : SELECT_OP
      generic map ( num_inputs => 6, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => X_Logic0_port, 
         -- Connections to port 'DATA3'
         DATA(2) => X_Logic0_port, 
         -- Connections to port 'DATA4'
         DATA(3) => X_Logic0_port, 
         -- Connections to port 'DATA5'
         DATA(4) => N526, 
         -- Connections to port 'DATA6'
         DATA(5) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N68, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N69, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N70, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N71, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N72, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N73, 
         -- Connections to port 'Z'
         Z(0) => key_en );
   C2123_cell : SELECT_OP
      generic map ( num_inputs => 6, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => X_Logic0_port, 
         -- Connections to port 'DATA3'
         DATA(2) => X_Logic0_port, 
         -- Connections to port 'DATA4'
         DATA(3) => X_Logic0_port, 
         -- Connections to port 'DATA5'
         DATA(4) => X_Logic0_port, 
         -- Connections to port 'DATA6'
         DATA(5) => N572, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N68, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N69, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N70, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N71, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N72, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N73, 
         -- Connections to port 'Z'
         Z(0) => msg_auth_valid_port );
   C2124_cell : SELECT_OP
      generic map ( num_inputs => 6, input_width => 4 )
      port map(
         -- Connections to port 'DATA1'
         DATA(3) => bdi_valid_bytes_3_port, DATA(2) => bdi_valid_bytes_2_port, 
               DATA(1) => bdi_valid_bytes_1_port, DATA(0) => 
               bdi_valid_bytes_0_port, 
         -- Connections to port 'DATA2'
         DATA(7) => bdi_valid_bytes_3_port, DATA(6) => bdi_valid_bytes_2_port, 
               DATA(5) => bdi_valid_bytes_1_port, DATA(4) => 
               bdi_valid_bytes_0_port, 
         -- Connections to port 'DATA3'
         DATA(11) => bdi_valid_bytes_3_port, DATA(10) => bdi_valid_bytes_2_port
               , DATA(9) => bdi_valid_bytes_1_port, DATA(8) => 
               bdi_valid_bytes_0_port, 
         -- Connections to port 'DATA4'
         DATA(15) => bdi_valid_bytes_3_port, DATA(14) => bdi_valid_bytes_2_port
               , DATA(13) => bdi_valid_bytes_1_port, DATA(12) => 
               bdi_valid_bytes_0_port, 
         -- Connections to port 'DATA5'
         DATA(19) => bdi_valid_bytes_3_port, DATA(18) => bdi_valid_bytes_2_port
               , DATA(17) => bdi_valid_bytes_1_port, DATA(16) => 
               bdi_valid_bytes_0_port, 
         -- Connections to port 'DATA6'
         DATA(23) => N562, DATA(22) => N561, DATA(21) => N560, DATA(20) => N559
               , 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N68, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N69, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N70, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N71, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N72, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N73, 
         -- Connections to port 'Z'
         Z(3) => bdo_valid_bytes_3_port, Z(2) => bdo_valid_bytes_2_port, Z(1) 
               => bdo_valid_bytes_1_port, Z(0) => bdo_valid_bytes_0_port );
   C2125_cell : SELECT_OP
      generic map ( num_inputs => 6, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => X_Logic0_port, 
         -- Connections to port 'DATA3'
         DATA(2) => X_Logic0_port, 
         -- Connections to port 'DATA4'
         DATA(3) => X_Logic0_port, 
         -- Connections to port 'DATA5'
         DATA(4) => X_Logic0_port, 
         -- Connections to port 'DATA6'
         DATA(5) => N569, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N68, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N69, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N70, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N71, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N72, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N73, 
         -- Connections to port 'Z'
         Z(0) => msg_auth_port );
   C2126_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 3 )
      port map(
         -- Connections to port 'DATA1'
         DATA(2) => X_Logic0_port, DATA(1) => X_Logic0_port, DATA(0) => 
               X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(5) => n_cyc_s_2_port, DATA(4) => n_cyc_s_1_port, DATA(3) => 
               n_cyc_s_0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N74, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N75, 
         -- Connections to port 'Z'
         Z(2) => N576, Z(1) => N575, Z(0) => N574 );
   B_74 : GTECH_BUF port map( A => rst, Z => N74);
   B_75 : GTECH_BUF port map( A => N573, Z => N75);
   C2127_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic1_port, 
         -- Connections to port 'DATA2'
         DATA(1) => hash_in_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N74, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N75, 
         -- Connections to port 'Z'
         Z(0) => N577 );
   C2128_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => n_tag_verified, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N74, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N75, 
         -- Connections to port 'Z'
         Z(0) => N578 );
   C2129_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 3 )
      port map(
         -- Connections to port 'DATA1'
         DATA(2) => X_Logic0_port, DATA(1) => X_Logic0_port, DATA(0) => 
               X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(5) => n_calling_state_2_port, DATA(4) => n_calling_state_1_port, 
               DATA(3) => n_calling_state_0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N74, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N75, 
         -- Connections to port 'Z'
         Z(2) => N581, Z(1) => N580, Z(0) => N579 );
   C2130_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => n_gtr_one_perm, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N74, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N75, 
         -- Connections to port 'Z'
         Z(0) => N582 );
   C2131_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => n_decrypt_op_s, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N74, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N75, 
         -- Connections to port 'Z'
         Z(0) => N583 );
   C2132_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => n_bdi_eot_prev, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N74, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N75, 
         -- Connections to port 'Z'
         Z(0) => N584 );
         X_Logic1_port <= '1';
         X_Logic0_port <= '0';
   B_76 : GTECH_BUF port map( A => N758, Z => xor_sel);
   I_69 : GTECH_NOT port map( A => cyc_s_2_port, Z => N76);
   I_70 : GTECH_NOT port map( A => N80, Z => N81);
   I_71 : GTECH_NOT port map( A => N83, Z => N84);
   I_72 : GTECH_NOT port map( A => N86, Z => N87);
   I_73 : GTECH_NOT port map( A => N89, Z => N90);
   I_74 : GTECH_NOT port map( A => N92, Z => N93);
   B_77 : GTECH_BUF port map( A => N78, Z => state_main_sel_5_port);
   C2160 : GTECH_OR2 port map( A => key_valid_port, B => bdi_valid_port, Z => 
                           N94);
   I_75 : GTECH_NOT port map( A => N94, Z => N95);
   I_76 : GTECH_NOT port map( A => hash_in_port, Z => N96);
   I_77 : GTECH_NOT port map( A => key_update_port, Z => N97);
   I_78 : GTECH_NOT port map( A => key_valid_port, Z => N102);
   B_78 : GTECH_BUF port map( A => N84, Z => N174);
   I_79 : GTECH_NOT port map( A => bdi_valid_port, Z => N175);
   C2182 : GTECH_AND2 port map( A => N174, B => N749, Z => N182);
   C2183 : GTECH_AND2 port map( A => N747, B => bdi_eot_port, Z => N183);
   I_80 : GTECH_NOT port map( A => N183, Z => N184);
   C2186 : GTECH_AND2 port map( A => N182, B => N184, Z => N185);
   C2187 : GTECH_OR2 port map( A => N734, B => N737, Z => N186);
   I_81 : GTECH_NOT port map( A => N186, Z => N187);
   C2190 : GTECH_AND2 port map( A => N185, B => N186, Z => N188);
   C2191 : GTECH_OR2 port map( A => N802, B => N728, Z => N189);
   C2192 : GTECH_OR2 port map( A => N722, B => N724, Z => N802);
   I_82 : GTECH_NOT port map( A => N189, Z => N190);
   C2195 : GTECH_AND2 port map( A => N188, B => N189, Z => N191);
   C2196 : GTECH_AND2 port map( A => N191, B => bdi_valid_port, Z => N192);
   C2200 : GTECH_AND2 port map( A => N192, B => bdi_eot_port, Z => N193);
   I_83 : GTECH_NOT port map( A => N657, Z => N194);
   C2203 : GTECH_AND2 port map( A => N193, B => N657, Z => N195);
   I_84 : GTECH_NOT port map( A => N196, Z => N197);
   C2206 : GTECH_AND2 port map( A => N195, B => N197, Z => n_1168);
   C2208 : GTECH_AND2 port map( A => N192, B => N752, Z => N205);
   C2209 : GTECH_AND2 port map( A => N712, B => N715, Z => N206);
   I_85 : GTECH_NOT port map( A => N206, Z => N207);
   C2212 : GTECH_AND2 port map( A => N696, B => N699, Z => N208);
   I_86 : GTECH_NOT port map( A => N208, Z => N209);
   I_87 : GTECH_NOT port map( A => N216, Z => N217);
   C2217 : GTECH_AND2 port map( A => N205, B => N217, Z => n_1169);
   C2219 : GTECH_AND2 port map( A => N724, B => N657, Z => N229);
   I_88 : GTECH_NOT port map( A => N229, Z => N230);
   C2222 : GTECH_AND2 port map( A => N185, B => N187, Z => N248);
   C2224 : GTECH_OR2 port map( A => N803, B => N724, Z => N249);
   C2225 : GTECH_OR2 port map( A => N640, B => N624, Z => N803);
   I_89 : GTECH_NOT port map( A => N249, Z => N250);
   C2228 : GTECH_AND2 port map( A => N248, B => N249, Z => N251);
   C2229 : GTECH_AND2 port map( A => bdi_valid_port, B => bdo_ready_port, Z => 
                           N252);
   I_90 : GTECH_NOT port map( A => N252, Z => N253);
   C2232 : GTECH_AND2 port map( A => N251, B => N252, Z => N254);
   C2233 : GTECH_AND2 port map( A => N254, B => bdi_eot_port, Z => N255);
   C2236 : GTECH_AND2 port map( A => N255, B => N661, Z => n_1170);
   C2238 : GTECH_AND2 port map( A => N254, B => N752, Z => n_1171);
   B_79 : GTECH_BUF port map( A => N87, Z => N317);
   C2243 : GTECH_AND2 port map( A => N805, B => N747, Z => N318);
   C2244 : GTECH_AND2 port map( A => N804, B => N752, Z => N805);
   C2245 : GTECH_AND2 port map( A => N724, B => N751, Z => N804);
   I_91 : GTECH_NOT port map( A => N318, Z => N319);
   C2248 : GTECH_AND2 port map( A => N317, B => N319, Z => N320);
   C2251 : GTECH_AND2 port map( A => N320, B => N742, Z => N321);
   C2254 : GTECH_AND2 port map( A => N321, B => N740, Z => N322);
   I_92 : GTECH_NOT port map( A => N323, Z => N324);
   C2257 : GTECH_AND2 port map( A => N322, B => N324, Z => n_1172);
   C2262 : GTECH_AND2 port map( A => N322, B => N722, Z => n_1173);
   C2263 : GTECH_AND2 port map( A => N806, B => N329, Z => N330);
   C2264 : GTECH_AND2 port map( A => bdi_valid_port, B => N707, Z => N806);
   I_93 : GTECH_NOT port map( A => N330, Z => N331);
   C2271 : GTECH_AND2 port map( A => N321, B => N739, Z => N356);
   C2274 : GTECH_AND2 port map( A => N356, B => N731, Z => N357);
   C2275 : GTECH_AND2 port map( A => N639, B => N623, Z => N358);
   I_94 : GTECH_NOT port map( A => N358, Z => N359);
   C2278 : GTECH_AND2 port map( A => N357, B => N358, Z => n_1174);
   C2280 : GTECH_AND2 port map( A => N357, B => N359, Z => N362);
   C2281 : GTECH_AND2 port map( A => N808, B => N363, Z => N364);
   C2282 : GTECH_AND2 port map( A => N807, B => N707, Z => N808);
   C2283 : GTECH_AND2 port map( A => bdi_valid_port, B => bdo_ready_port, Z => 
                           N807);
   I_95 : GTECH_NOT port map( A => N364, Z => N365);
   C2286 : GTECH_AND2 port map( A => N362, B => N364, Z => N366);
   C2288 : GTECH_AND2 port map( A => N366, B => bdi_eot_port, Z => n_1175);
   C2290 : GTECH_AND2 port map( A => N366, B => N752, Z => n_1176);
   C2301 : GTECH_AND2 port map( A => bdi_valid_port, B => N692, Z => N408);
   I_96 : GTECH_NOT port map( A => N408, Z => N409);
   C2307 : GTECH_OR2 port map( A => N686, B => N689, Z => N510);
   I_97 : GTECH_NOT port map( A => N510, Z => N511);
   B_80 : GTECH_BUF port map( A => N93, Z => N527);
   C2318 : GTECH_AND2 port map( A => N652, B => N654, Z => N528);
   I_98 : GTECH_NOT port map( A => N528, Z => N529);
   C2321 : GTECH_AND2 port map( A => N527, B => decrypt_op_s, Z => N542);
   C2322 : GTECH_AND2 port map( A => bdi_valid_port, B => msg_auth_ready, Z => 
                           N543);
   I_99 : GTECH_NOT port map( A => N543, Z => N544);
   C2325 : GTECH_AND2 port map( A => N542, B => N543, Z => N545);
   C2328 : GTECH_AND2 port map( A => N545, B => N682, Z => n_1177);
   I_100 : GTECH_NOT port map( A => N546, Z => N547);
   C2331 : GTECH_AND2 port map( A => N545, B => N681, Z => n_1178);
   I_101 : GTECH_NOT port map( A => rst, Z => N573);
   C2336 : GTECH_AND2 port map( A => state_main_sel_5_port, B => N573, Z => 
                           N585);
   C2337 : GTECH_AND2 port map( A => N95, B => N585, Z => N586);
   C2338 : GTECH_AND2 port map( A => N81, B => N573, Z => N587);
   C2339 : GTECH_AND2 port map( A => key_valid_port, B => N587, Z => N588);
   C2340 : GTECH_OR2 port map( A => N586, B => N588, Z => N589);
   C2341 : GTECH_AND2 port map( A => N93, B => N573, Z => N590);
   C2342 : GTECH_AND2 port map( A => decrypt_op_s, B => N590, Z => N591);
   C2343 : GTECH_AND2 port map( A => N544, B => N591, Z => N592);
   C2344 : GTECH_OR2 port map( A => N589, B => N592, Z => N593);
   I_102 : GTECH_NOT port map( A => N593, Z => N594);
   C2346 : GTECH_OR2 port map( A => N586, B => N587, Z => N595);
   C2347 : GTECH_AND2 port map( A => N84, B => N573, Z => N596);
   C2348 : GTECH_OR2 port map( A => N595, B => N596, Z => N597);
   C2349 : GTECH_AND2 port map( A => N87, B => N573, Z => N598);
   C2350 : GTECH_OR2 port map( A => N597, B => N598, Z => N599);
   C2351 : GTECH_AND2 port map( A => N90, B => N573, Z => N600);
   C2352 : GTECH_OR2 port map( A => N599, B => N600, Z => N601);
   C2353 : GTECH_OR2 port map( A => N601, B => N590, Z => N602);
   I_103 : GTECH_NOT port map( A => N602, Z => N603);
   C2355 : GTECH_AND2 port map( A => N94, B => N585, Z => N604);
   C2356 : GTECH_AND2 port map( A => N96, B => N604, Z => N605);
   C2357 : GTECH_AND2 port map( A => key_update_port, B => N605, Z => N606);
   C2358 : GTECH_OR2 port map( A => N606, B => N586, Z => N607);
   C2359 : GTECH_OR2 port map( A => N607, B => N588, Z => N608);
   C2360 : GTECH_OR2 port map( A => N608, B => N596, Z => N609);
   C2361 : GTECH_OR2 port map( A => N609, B => N591, Z => N610);
   I_104 : GTECH_NOT port map( A => N610, Z => N611);
   C2363 : GTECH_OR2 port map( A => N587, B => N596, Z => N612);
   C2364 : GTECH_OR2 port map( A => N612, B => N600, Z => N613);
   C2365 : GTECH_OR2 port map( A => N613, B => N590, Z => N614);
   I_105 : GTECH_NOT port map( A => N614, Z => N615);
   C2367 : GTECH_OR2 port map( A => N605, B => N586, Z => N616);
   C2368 : GTECH_OR2 port map( A => N616, B => N587, Z => N617);
   C2369 : GTECH_OR2 port map( A => N617, B => N598, Z => N618);
   C2370 : GTECH_OR2 port map( A => N618, B => N600, Z => N619);
   C2371 : GTECH_OR2 port map( A => N619, B => N590, Z => N620);
   I_106 : GTECH_NOT port map( A => N620, Z => N621);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_LWC_1.all;

entity PreProcessor_2 is

   port( clk, rst : in std_logic;  pdi_data : in std_logic_vector (31 downto 0)
         ;  pdi_valid : in std_logic;  pdi_ready : out std_logic;  sdi_data : 
         in std_logic_vector (31 downto 0);  sdi_valid : in std_logic;  
         sdi_ready : out std_logic;  key : out std_logic_vector (31 downto 0); 
         key_valid : out std_logic;  key_ready : in std_logic;  bdi : out 
         std_logic_vector (31 downto 0);  bdi_valid : out std_logic;  bdi_ready
         : in std_logic;  bdi_pad_loc, bdi_valid_bytes : out std_logic_vector 
         (3 downto 0);  bdi_size : out std_logic_vector (2 downto 0);  bdi_eot,
         bdi_eoi : out std_logic;  bdi_type : out std_logic_vector (3 downto 0)
         ;  decrypt, hash, key_update : out std_logic;  cmd : out 
         std_logic_vector (31 downto 0);  cmd_valid : out std_logic;  cmd_ready
         : in std_logic);

end PreProcessor_2;

architecture SYN_PreProcessor of PreProcessor_2 is

   component GTECH_NOT
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component GTECH_OR2
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component GTECH_AND2
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component GTECH_BUF
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
      generic ( ac_as_q, ac_as_qn, sc_ss_q : integer );
      port(
         clear, preset, enable, data_in, synch_clear, synch_preset, 
            synch_toggle, synch_enable, next_state, clocked_on : in std_logic;
         Q, QN : buffer std_logic
      );
   end component;
   
   component DATA_PISO_2
      port( clk, rst : in std_logic;  data_size_p : in std_logic_vector (2 
            downto 0);  data_size_s : out std_logic_vector (2 downto 0);  
            data_s : out std_logic_vector (31 downto 0);  data_valid_s : out 
            std_logic;  data_ready_s : in std_logic;  data_p : in 
            std_logic_vector (31 downto 0);  data_valid_p : in std_logic;  
            data_ready_p : out std_logic;  valid_bytes_p : in std_logic_vector 
            (3 downto 0);  valid_bytes_s : out std_logic_vector (3 downto 0);  
            pad_loc_p : in std_logic_vector (3 downto 0);  pad_loc_s : out 
            std_logic_vector (3 downto 0);  eoi_p : in std_logic;  eoi_s : out 
            std_logic;  eot_p : in std_logic;  eot_s : out std_logic);
   end component;
   
   component KEY_PISO_2
      port( clk, rst : in std_logic;  data_s : out std_logic_vector (31 downto 
            0);  data_valid_s : out std_logic;  data_ready_s : in std_logic;  
            data_p : in std_logic_vector (31 downto 0);  data_valid_p : in 
            std_logic;  data_ready_p : out std_logic);
   end component;
   
   component StepDownCountLd_N16_step4_2
      port( clk, len, ena : in std_logic;  load : in std_logic_vector (15 
            downto 0);  count : out std_logic_vector (15 downto 0));
   end component;
   
   signal N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15,
      N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30
      , N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, 
      N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59
      , N60, N61, N62, N63, X_Logic1_port, X_Logic0_port, clk_port, 
      pdi_valid_port, pdi_ready_port, sdi_data_31_port, sdi_data_30_port, 
      sdi_data_29_port, sdi_data_28_port, sdi_data_27_port, sdi_data_26_port, 
      sdi_data_25_port, sdi_data_24_port, sdi_data_23_port, sdi_data_22_port, 
      sdi_data_21_port, sdi_data_20_port, sdi_data_19_port, sdi_data_18_port, 
      sdi_data_17_port, sdi_data_16_port, sdi_data_15_port, sdi_data_14_port, 
      sdi_data_13_port, sdi_data_12_port, sdi_data_11_port, sdi_data_10_port, 
      sdi_data_9_port, sdi_data_8_port, sdi_data_7_port, sdi_data_6_port, 
      sdi_data_5_port, sdi_data_4_port, sdi_data_3_port, sdi_data_2_port, 
      sdi_data_1_port, sdi_data_0_port, sdi_valid_port, sdi_ready_port, 
      bdi_type_3_port, bdi_type_2_port, bdi_type_1_port, bdi_type_0_port, 
      decrypt_port, hash_port, key_update_port, cmd_31_port, cmd_30_port, 
      cmd_29_port, cmd_28_port, cmd_27_port, cmd_26_port, cmd_25_port, 
      cmd_24_port, cmd_23_port, cmd_22_port, cmd_21_port, cmd_20_port, 
      cmd_19_port, cmd_18_port, cmd_17_port, cmd_16_port, cmd_15_port, 
      cmd_14_port, cmd_13_port, cmd_12_port, cmd_11_port, cmd_10_port, 
      cmd_9_port, cmd_8_port, cmd_7_port, cmd_6_port, cmd_5_port, cmd_4_port, 
      cmd_3_port, cmd_2_port, cmd_1_port, cmd_0_port, cmd_valid_port, 
      cmd_ready_port, len_SegLenCnt, en_SegLenCnt, load_SegLenCnt_15_port, 
      load_SegLenCnt_14_port, load_SegLenCnt_13_port, load_SegLenCnt_12_port, 
      load_SegLenCnt_11_port, load_SegLenCnt_10_port, load_SegLenCnt_9_port, 
      load_SegLenCnt_8_port, load_SegLenCnt_7_port, load_SegLenCnt_6_port, 
      load_SegLenCnt_5_port, load_SegLenCnt_4_port, load_SegLenCnt_3_port, 
      load_SegLenCnt_2_port, load_SegLenCnt_1_port, load_SegLenCnt_0_port, 
      dout_SegLenCnt_15_port, dout_SegLenCnt_14_port, dout_SegLenCnt_13_port, 
      dout_SegLenCnt_12_port, dout_SegLenCnt_11_port, dout_SegLenCnt_10_port, 
      dout_SegLenCnt_9_port, dout_SegLenCnt_8_port, dout_SegLenCnt_7_port, 
      dout_SegLenCnt_6_port, dout_SegLenCnt_5_port, dout_SegLenCnt_4_port, 
      dout_SegLenCnt_3_port, dout_SegLenCnt_2_port, dout_SegLenCnt_1_port, 
      dout_SegLenCnt_0_port, N64, last_flit_of_segment, N65, N66, N67, N68, N69
      , N70, N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, 
      N84, N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98
      , N99, N100, N101, N102, N103, N104, N105, N106, N107, N108, N109, N110, 
      N111, N112, N113, N114, N115, N116, N117, N118, N119, N120, N121, N122, 
      N123, N124, N125, N126, N127, N128, N129, N130, N131, N132, N133, N134, 
      bdi_valid_bytes_p_3_port, bdi_valid_bytes_p_2_port, 
      bdi_valid_bytes_p_1_port, bdi_valid_bytes_p_0_port, N135, N136, N137, 
      N138, N139, N140, N141, N142, N143, N144, N145, N146, N147, N148, N149, 
      N150, N151, N152, N153, N154, N155, N156, N157, N158, N159, N160, N161, 
      N162, N163, N164, N165, N166, N167, N168, N169, N170, N171, N172, N173, 
      N174, N175, N176, N177, N178, N179, N180, N181, N182, N183, N184, N185, 
      N186, N187, N188, N189, N190, N191, N192, N193, N194, N195, N196, N197, 
      N198, N199, N200, N201, N202, bdi_pad_loc_p_3_port, bdi_pad_loc_p_2_port,
      bdi_pad_loc_p_1_port, bdi_pad_loc_p_0_port, eoi_flag, eot_flag, 
      sel_sdi_length, N203, N204, bdi_size_p_2_port, bdi_size_p_1_port, 
      bdi_size_p_0_port, bdi_eoi_internal, bdi_eot_internal, key_ready_p, 
      key_valid_p, bdi_ready_p, bdi_valid_p, N205, pr_state_3_port, 
      pr_state_2_port, pr_state_1_port, pr_state_0_port, nx_state_3_port, 
      nx_state_2_port, nx_state_1_port, nx_state_0_port, N206, N207, N208, N209
      , N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220, N221,
      N222, N223, N224, N225, N226, N227, N228, N229, N230, N231, N232, N233, 
      N234, N235, N236, N237, N238, N239, N240, N241, N242, N243, N244, N245, 
      N246, N247, N248, N249, N250, N251, N252, N253, N254, N255, N256, N257, 
      N258, N259, N260, N261, N262, N263, N264, N265, N266, N267, N268, N269, 
      N270, N271, N272, N273, N274, N275, N276, N277, N278, N279, N280, N281, 
      N282, N283, N284, N285, N286, N287, N288, N289, N290, N291, N292, N293, 
      N294, N295, N296, N297, N298, N299, N300, N301, N302, N303, N304, N305, 
      N306, N307, N308, N309, N310, N311, N312, N313, N314, N315, N316, N317, 
      N318, N319, N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, 
      N330, N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341, 
      N342, N343, N344, N345, N346, N347, N348, N349, N350, N351, N352, N353, 
      N354, N355, N356, N357, N358, N359, N360, N361, N362, N363, N364, N365, 
      N366, N367, N368, N369, N370, N371, N372, N373, N374, N375, N376, N377, 
      N378, N379, N380, N381, N382, N383, N384, N385, N386, N387, N388, N389, 
      N390, N391, N392, N393, N394, N395, N396, N397, N398, N399, N400, N401, 
      N402, N403, N404, N405, N406, N407, N408, N409, N410, N411, N412, N413, 
      N414, N415, N416, N417, N418, N419, N420, N421, N422, N423, N424, N425, 
      N426, N427, N428, N429, N430, N431, N432, N433, N434, N435, N436, N437, 
      N438, N439, N440, N441, N442, N443, N444, N445, N446, N447, N448, N449, 
      N450, N451, N452, N453, N454, N455, N456, N457, N458, N459, N460, N461, 
      N462, N463, N464, N465, N466, N467, N468, N469, N470, N471, N472, N473, 
      N474, N475, N476, N477, N478, N479, N480, N481, N482, N483, N484, N485, 
      N486, N487, N488, N489, N490, N491, N492, N493, N494, N495, N496, N497, 
      N498, N499, N500, N501, N502, N503, N504, N505, N506, N507, N508, N509, 
      N510, N511, N512, N513, N514, N515, N516, N517, N518, N519, N520, N521, 
      N522, N523, N524, N525, N526, N527, N528, N529, N530, N531, N532, n_1179,
      n_1180, n_1181, n_1182, n_1183, n_1184, n_1185, n_1186 : std_logic;

begin
   clk_port <= clk;
   ( cmd_31_port, cmd_30_port, cmd_29_port, cmd_28_port, cmd_27_port, 
      cmd_26_port, cmd_25_port, cmd_24_port, cmd_23_port, cmd_22_port, 
      cmd_21_port, cmd_20_port, cmd_19_port, cmd_18_port, cmd_17_port, 
      cmd_16_port, cmd_15_port, cmd_14_port, cmd_13_port, cmd_12_port, 
      cmd_11_port, cmd_10_port, cmd_9_port, cmd_8_port, cmd_7_port, cmd_6_port,
      cmd_5_port, cmd_4_port, cmd_3_port, cmd_2_port, cmd_1_port, cmd_0_port ) 
      <= pdi_data;
   pdi_valid_port <= pdi_valid;
   pdi_ready <= pdi_ready_port;
   ( sdi_data_31_port, sdi_data_30_port, sdi_data_29_port, sdi_data_28_port, 
      sdi_data_27_port, sdi_data_26_port, sdi_data_25_port, sdi_data_24_port, 
      sdi_data_23_port, sdi_data_22_port, sdi_data_21_port, sdi_data_20_port, 
      sdi_data_19_port, sdi_data_18_port, sdi_data_17_port, sdi_data_16_port, 
      sdi_data_15_port, sdi_data_14_port, sdi_data_13_port, sdi_data_12_port, 
      sdi_data_11_port, sdi_data_10_port, sdi_data_9_port, sdi_data_8_port, 
      sdi_data_7_port, sdi_data_6_port, sdi_data_5_port, sdi_data_4_port, 
      sdi_data_3_port, sdi_data_2_port, sdi_data_1_port, sdi_data_0_port ) <= 
      sdi_data;
   sdi_valid_port <= sdi_valid;
   sdi_ready <= sdi_ready_port;
   bdi_type <= ( bdi_type_3_port, bdi_type_2_port, bdi_type_1_port, 
      bdi_type_0_port );
   decrypt <= decrypt_port;
   hash <= hash_port;
   key_update <= key_update_port;
   cmd <= ( cmd_31_port, cmd_30_port, cmd_29_port, cmd_28_port, cmd_27_port, 
      cmd_26_port, cmd_25_port, cmd_24_port, cmd_23_port, cmd_22_port, 
      cmd_21_port, cmd_20_port, cmd_19_port, cmd_18_port, cmd_17_port, 
      cmd_16_port, cmd_15_port, cmd_14_port, cmd_13_port, cmd_12_port, 
      cmd_11_port, cmd_10_port, cmd_9_port, cmd_8_port, cmd_7_port, cmd_6_port,
      cmd_5_port, cmd_4_port, cmd_3_port, cmd_2_port, cmd_1_port, cmd_0_port );
   cmd_valid <= cmd_valid_port;
   cmd_ready_port <= cmd_ready;
   
   SegLen : StepDownCountLd_N16_step4_2 port map( clk => clk_port, len => 
                           len_SegLenCnt, ena => en_SegLenCnt, load(15) => 
                           load_SegLenCnt_15_port, load(14) => 
                           load_SegLenCnt_14_port, load(13) => 
                           load_SegLenCnt_13_port, load(12) => 
                           load_SegLenCnt_12_port, load(11) => 
                           load_SegLenCnt_11_port, load(10) => 
                           load_SegLenCnt_10_port, load(9) => 
                           load_SegLenCnt_9_port, load(8) => 
                           load_SegLenCnt_8_port, load(7) => 
                           load_SegLenCnt_7_port, load(6) => 
                           load_SegLenCnt_6_port, load(5) => 
                           load_SegLenCnt_5_port, load(4) => 
                           load_SegLenCnt_4_port, load(3) => 
                           load_SegLenCnt_3_port, load(2) => 
                           load_SegLenCnt_2_port, load(1) => 
                           load_SegLenCnt_1_port, load(0) => 
                           load_SegLenCnt_0_port, count(15) => 
                           dout_SegLenCnt_15_port, count(14) => 
                           dout_SegLenCnt_14_port, count(13) => 
                           dout_SegLenCnt_13_port, count(12) => 
                           dout_SegLenCnt_12_port, count(11) => 
                           dout_SegLenCnt_11_port, count(10) => 
                           dout_SegLenCnt_10_port, count(9) => 
                           dout_SegLenCnt_9_port, count(8) => 
                           dout_SegLenCnt_8_port, count(7) => 
                           dout_SegLenCnt_7_port, count(6) => 
                           dout_SegLenCnt_6_port, count(5) => 
                           dout_SegLenCnt_5_port, count(4) => 
                           dout_SegLenCnt_4_port, count(3) => 
                           dout_SegLenCnt_3_port, count(2) => 
                           dout_SegLenCnt_2_port, count(1) => 
                           dout_SegLenCnt_1_port, count(0) => 
                           dout_SegLenCnt_0_port);
   lte_155 : process ( dout_SegLenCnt_15_port, dout_SegLenCnt_14_port, 
         dout_SegLenCnt_13_port, dout_SegLenCnt_12_port, dout_SegLenCnt_11_port
         , dout_SegLenCnt_10_port, dout_SegLenCnt_9_port, dout_SegLenCnt_8_port
         , dout_SegLenCnt_7_port, dout_SegLenCnt_6_port, dout_SegLenCnt_5_port,
         dout_SegLenCnt_4_port, dout_SegLenCnt_3_port, dout_SegLenCnt_2_port, 
         dout_SegLenCnt_1_port, dout_SegLenCnt_0_port, X_Logic0_port, 
         X_Logic1_port )
      variable A : UNSIGNED( 15 downto 0 );
      variable B : UNSIGNED( 15 downto 0 );
      variable Z : UNSIGNED( 0 downto 0 );
   begin
      A := ( dout_SegLenCnt_15_port, dout_SegLenCnt_14_port, 
            dout_SegLenCnt_13_port, dout_SegLenCnt_12_port, 
            dout_SegLenCnt_11_port, dout_SegLenCnt_10_port, 
            dout_SegLenCnt_9_port, dout_SegLenCnt_8_port, dout_SegLenCnt_7_port
            , dout_SegLenCnt_6_port, dout_SegLenCnt_5_port, 
            dout_SegLenCnt_4_port, dout_SegLenCnt_3_port, dout_SegLenCnt_2_port
            , dout_SegLenCnt_1_port, dout_SegLenCnt_0_port );
      B := ( X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
            X_Logic0_port, X_Logic1_port, X_Logic0_port, X_Logic0_port );
      if ( A <= B ) then
         Z := ( others => '1' );
      else
         Z := ( others => '0' );
      end if;
      ( 0 => N64 ) <= Z;
   end process;
   
   C14 : GTECH_OR2 port map( A => dout_SegLenCnt_14_port, B => 
                           dout_SegLenCnt_15_port, Z => N65);
   C15 : GTECH_OR2 port map( A => dout_SegLenCnt_13_port, B => N65, Z => N66);
   C16 : GTECH_OR2 port map( A => dout_SegLenCnt_12_port, B => N66, Z => N67);
   C17 : GTECH_OR2 port map( A => dout_SegLenCnt_11_port, B => N67, Z => N68);
   C18 : GTECH_OR2 port map( A => dout_SegLenCnt_10_port, B => N68, Z => N69);
   C19 : GTECH_OR2 port map( A => dout_SegLenCnt_9_port, B => N69, Z => N70);
   C20 : GTECH_OR2 port map( A => dout_SegLenCnt_8_port, B => N70, Z => N71);
   C21 : GTECH_OR2 port map( A => dout_SegLenCnt_7_port, B => N71, Z => N72);
   C22 : GTECH_OR2 port map( A => dout_SegLenCnt_6_port, B => N72, Z => N73);
   C23 : GTECH_OR2 port map( A => dout_SegLenCnt_5_port, B => N73, Z => N74);
   C24 : GTECH_OR2 port map( A => dout_SegLenCnt_4_port, B => N74, Z => N75);
   C25 : GTECH_OR2 port map( A => dout_SegLenCnt_3_port, B => N75, Z => N76);
   C26 : GTECH_OR2 port map( A => dout_SegLenCnt_2_port, B => N76, Z => N77);
   C27 : GTECH_OR2 port map( A => dout_SegLenCnt_1_port, B => N77, Z => N78);
   C28 : GTECH_OR2 port map( A => dout_SegLenCnt_0_port, B => N78, Z => N79);
   I_0 : GTECH_NOT port map( A => N79, Z => N80);
   I_1 : GTECH_NOT port map( A => dout_SegLenCnt_0_port, Z => N81);
   C31 : GTECH_OR2 port map( A => dout_SegLenCnt_14_port, B => 
                           dout_SegLenCnt_15_port, Z => N82);
   C32 : GTECH_OR2 port map( A => dout_SegLenCnt_13_port, B => N82, Z => N83);
   C33 : GTECH_OR2 port map( A => dout_SegLenCnt_12_port, B => N83, Z => N84);
   C34 : GTECH_OR2 port map( A => dout_SegLenCnt_11_port, B => N84, Z => N85);
   C35 : GTECH_OR2 port map( A => dout_SegLenCnt_10_port, B => N85, Z => N86);
   C36 : GTECH_OR2 port map( A => dout_SegLenCnt_9_port, B => N86, Z => N87);
   C37 : GTECH_OR2 port map( A => dout_SegLenCnt_8_port, B => N87, Z => N88);
   C38 : GTECH_OR2 port map( A => dout_SegLenCnt_7_port, B => N88, Z => N89);
   C39 : GTECH_OR2 port map( A => dout_SegLenCnt_6_port, B => N89, Z => N90);
   C40 : GTECH_OR2 port map( A => dout_SegLenCnt_5_port, B => N90, Z => N91);
   C41 : GTECH_OR2 port map( A => dout_SegLenCnt_4_port, B => N91, Z => N92);
   C42 : GTECH_OR2 port map( A => dout_SegLenCnt_3_port, B => N92, Z => N93);
   C43 : GTECH_OR2 port map( A => dout_SegLenCnt_2_port, B => N93, Z => N94);
   C44 : GTECH_OR2 port map( A => dout_SegLenCnt_1_port, B => N94, Z => N95);
   C45 : GTECH_OR2 port map( A => N81, B => N95, Z => N96);
   I_2 : GTECH_NOT port map( A => N96, Z => N97);
   I_3 : GTECH_NOT port map( A => dout_SegLenCnt_1_port, Z => N98);
   C48 : GTECH_OR2 port map( A => dout_SegLenCnt_14_port, B => 
                           dout_SegLenCnt_15_port, Z => N99);
   C49 : GTECH_OR2 port map( A => dout_SegLenCnt_13_port, B => N99, Z => N100);
   C50 : GTECH_OR2 port map( A => dout_SegLenCnt_12_port, B => N100, Z => N101)
                           ;
   C51 : GTECH_OR2 port map( A => dout_SegLenCnt_11_port, B => N101, Z => N102)
                           ;
   C52 : GTECH_OR2 port map( A => dout_SegLenCnt_10_port, B => N102, Z => N103)
                           ;
   C53 : GTECH_OR2 port map( A => dout_SegLenCnt_9_port, B => N103, Z => N104);
   C54 : GTECH_OR2 port map( A => dout_SegLenCnt_8_port, B => N104, Z => N105);
   C55 : GTECH_OR2 port map( A => dout_SegLenCnt_7_port, B => N105, Z => N106);
   C56 : GTECH_OR2 port map( A => dout_SegLenCnt_6_port, B => N106, Z => N107);
   C57 : GTECH_OR2 port map( A => dout_SegLenCnt_5_port, B => N107, Z => N108);
   C58 : GTECH_OR2 port map( A => dout_SegLenCnt_4_port, B => N108, Z => N109);
   C59 : GTECH_OR2 port map( A => dout_SegLenCnt_3_port, B => N109, Z => N110);
   C60 : GTECH_OR2 port map( A => dout_SegLenCnt_2_port, B => N110, Z => N111);
   C61 : GTECH_OR2 port map( A => N98, B => N111, Z => N112);
   C62 : GTECH_OR2 port map( A => dout_SegLenCnt_0_port, B => N112, Z => N113);
   I_4 : GTECH_NOT port map( A => N113, Z => N114);
   C66 : GTECH_OR2 port map( A => dout_SegLenCnt_14_port, B => 
                           dout_SegLenCnt_15_port, Z => N115);
   C67 : GTECH_OR2 port map( A => dout_SegLenCnt_13_port, B => N115, Z => N116)
                           ;
   C68 : GTECH_OR2 port map( A => dout_SegLenCnt_12_port, B => N116, Z => N117)
                           ;
   C69 : GTECH_OR2 port map( A => dout_SegLenCnt_11_port, B => N117, Z => N118)
                           ;
   C70 : GTECH_OR2 port map( A => dout_SegLenCnt_10_port, B => N118, Z => N119)
                           ;
   C71 : GTECH_OR2 port map( A => dout_SegLenCnt_9_port, B => N119, Z => N120);
   C72 : GTECH_OR2 port map( A => dout_SegLenCnt_8_port, B => N120, Z => N121);
   C73 : GTECH_OR2 port map( A => dout_SegLenCnt_7_port, B => N121, Z => N122);
   C74 : GTECH_OR2 port map( A => dout_SegLenCnt_6_port, B => N122, Z => N123);
   C75 : GTECH_OR2 port map( A => dout_SegLenCnt_5_port, B => N123, Z => N124);
   C76 : GTECH_OR2 port map( A => dout_SegLenCnt_4_port, B => N124, Z => N125);
   C77 : GTECH_OR2 port map( A => dout_SegLenCnt_3_port, B => N125, Z => N126);
   C78 : GTECH_OR2 port map( A => dout_SegLenCnt_2_port, B => N126, Z => N127);
   C79 : GTECH_OR2 port map( A => N98, B => N127, Z => N128);
   C80 : GTECH_OR2 port map( A => N81, B => N128, Z => N129);
   I_5 : GTECH_NOT port map( A => N129, Z => N130);
   C99 : GTECH_OR2 port map( A => dout_SegLenCnt_14_port, B => 
                           dout_SegLenCnt_15_port, Z => N135);
   C100 : GTECH_OR2 port map( A => dout_SegLenCnt_13_port, B => N135, Z => N136
                           );
   C101 : GTECH_OR2 port map( A => dout_SegLenCnt_12_port, B => N136, Z => N137
                           );
   C102 : GTECH_OR2 port map( A => dout_SegLenCnt_11_port, B => N137, Z => N138
                           );
   C103 : GTECH_OR2 port map( A => dout_SegLenCnt_10_port, B => N138, Z => N139
                           );
   C104 : GTECH_OR2 port map( A => dout_SegLenCnt_9_port, B => N139, Z => N140)
                           ;
   C105 : GTECH_OR2 port map( A => dout_SegLenCnt_8_port, B => N140, Z => N141)
                           ;
   C106 : GTECH_OR2 port map( A => dout_SegLenCnt_7_port, B => N141, Z => N142)
                           ;
   C107 : GTECH_OR2 port map( A => dout_SegLenCnt_6_port, B => N142, Z => N143)
                           ;
   C108 : GTECH_OR2 port map( A => dout_SegLenCnt_5_port, B => N143, Z => N144)
                           ;
   C109 : GTECH_OR2 port map( A => dout_SegLenCnt_4_port, B => N144, Z => N145)
                           ;
   C110 : GTECH_OR2 port map( A => dout_SegLenCnt_3_port, B => N145, Z => N146)
                           ;
   C111 : GTECH_OR2 port map( A => dout_SegLenCnt_2_port, B => N146, Z => N147)
                           ;
   C112 : GTECH_OR2 port map( A => dout_SegLenCnt_1_port, B => N147, Z => N148)
                           ;
   C113 : GTECH_OR2 port map( A => dout_SegLenCnt_0_port, B => N148, Z => N149)
                           ;
   I_6 : GTECH_NOT port map( A => N149, Z => N150);
   C116 : GTECH_OR2 port map( A => dout_SegLenCnt_14_port, B => 
                           dout_SegLenCnt_15_port, Z => N151);
   C117 : GTECH_OR2 port map( A => dout_SegLenCnt_13_port, B => N151, Z => N152
                           );
   C118 : GTECH_OR2 port map( A => dout_SegLenCnt_12_port, B => N152, Z => N153
                           );
   C119 : GTECH_OR2 port map( A => dout_SegLenCnt_11_port, B => N153, Z => N154
                           );
   C120 : GTECH_OR2 port map( A => dout_SegLenCnt_10_port, B => N154, Z => N155
                           );
   C121 : GTECH_OR2 port map( A => dout_SegLenCnt_9_port, B => N155, Z => N156)
                           ;
   C122 : GTECH_OR2 port map( A => dout_SegLenCnt_8_port, B => N156, Z => N157)
                           ;
   C123 : GTECH_OR2 port map( A => dout_SegLenCnt_7_port, B => N157, Z => N158)
                           ;
   C124 : GTECH_OR2 port map( A => dout_SegLenCnt_6_port, B => N158, Z => N159)
                           ;
   C125 : GTECH_OR2 port map( A => dout_SegLenCnt_5_port, B => N159, Z => N160)
                           ;
   C126 : GTECH_OR2 port map( A => dout_SegLenCnt_4_port, B => N160, Z => N161)
                           ;
   C127 : GTECH_OR2 port map( A => dout_SegLenCnt_3_port, B => N161, Z => N162)
                           ;
   C128 : GTECH_OR2 port map( A => dout_SegLenCnt_2_port, B => N162, Z => N163)
                           ;
   C129 : GTECH_OR2 port map( A => dout_SegLenCnt_1_port, B => N163, Z => N164)
                           ;
   C130 : GTECH_OR2 port map( A => N81, B => N164, Z => N165);
   I_7 : GTECH_NOT port map( A => N165, Z => N166);
   C133 : GTECH_OR2 port map( A => dout_SegLenCnt_14_port, B => 
                           dout_SegLenCnt_15_port, Z => N167);
   C134 : GTECH_OR2 port map( A => dout_SegLenCnt_13_port, B => N167, Z => N168
                           );
   C135 : GTECH_OR2 port map( A => dout_SegLenCnt_12_port, B => N168, Z => N169
                           );
   C136 : GTECH_OR2 port map( A => dout_SegLenCnt_11_port, B => N169, Z => N170
                           );
   C137 : GTECH_OR2 port map( A => dout_SegLenCnt_10_port, B => N170, Z => N171
                           );
   C138 : GTECH_OR2 port map( A => dout_SegLenCnt_9_port, B => N171, Z => N172)
                           ;
   C139 : GTECH_OR2 port map( A => dout_SegLenCnt_8_port, B => N172, Z => N173)
                           ;
   C140 : GTECH_OR2 port map( A => dout_SegLenCnt_7_port, B => N173, Z => N174)
                           ;
   C141 : GTECH_OR2 port map( A => dout_SegLenCnt_6_port, B => N174, Z => N175)
                           ;
   C142 : GTECH_OR2 port map( A => dout_SegLenCnt_5_port, B => N175, Z => N176)
                           ;
   C143 : GTECH_OR2 port map( A => dout_SegLenCnt_4_port, B => N176, Z => N177)
                           ;
   C144 : GTECH_OR2 port map( A => dout_SegLenCnt_3_port, B => N177, Z => N178)
                           ;
   C145 : GTECH_OR2 port map( A => dout_SegLenCnt_2_port, B => N178, Z => N179)
                           ;
   C146 : GTECH_OR2 port map( A => N98, B => N179, Z => N180);
   C147 : GTECH_OR2 port map( A => dout_SegLenCnt_0_port, B => N180, Z => N181)
                           ;
   I_8 : GTECH_NOT port map( A => N181, Z => N182);
   C151 : GTECH_OR2 port map( A => dout_SegLenCnt_14_port, B => 
                           dout_SegLenCnt_15_port, Z => N183);
   C152 : GTECH_OR2 port map( A => dout_SegLenCnt_13_port, B => N183, Z => N184
                           );
   C153 : GTECH_OR2 port map( A => dout_SegLenCnt_12_port, B => N184, Z => N185
                           );
   C154 : GTECH_OR2 port map( A => dout_SegLenCnt_11_port, B => N185, Z => N186
                           );
   C155 : GTECH_OR2 port map( A => dout_SegLenCnt_10_port, B => N186, Z => N187
                           );
   C156 : GTECH_OR2 port map( A => dout_SegLenCnt_9_port, B => N187, Z => N188)
                           ;
   C157 : GTECH_OR2 port map( A => dout_SegLenCnt_8_port, B => N188, Z => N189)
                           ;
   C158 : GTECH_OR2 port map( A => dout_SegLenCnt_7_port, B => N189, Z => N190)
                           ;
   C159 : GTECH_OR2 port map( A => dout_SegLenCnt_6_port, B => N190, Z => N191)
                           ;
   C160 : GTECH_OR2 port map( A => dout_SegLenCnt_5_port, B => N191, Z => N192)
                           ;
   C161 : GTECH_OR2 port map( A => dout_SegLenCnt_4_port, B => N192, Z => N193)
                           ;
   C162 : GTECH_OR2 port map( A => dout_SegLenCnt_3_port, B => N193, Z => N194)
                           ;
   C163 : GTECH_OR2 port map( A => dout_SegLenCnt_2_port, B => N194, Z => N195)
                           ;
   C164 : GTECH_OR2 port map( A => N98, B => N195, Z => N196);
   C165 : GTECH_OR2 port map( A => N81, B => N196, Z => N197);
   I_9 : GTECH_NOT port map( A => N197, Z => N198);
   hash_internal_reg : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N426, next_state => N401, 
               clocked_on => clk_port, Q => hash_port, QN => n_1179);
   decrypt_internal_reg : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N426, next_state => N399, 
               clocked_on => clk_port, Q => decrypt_port, QN => n_1180);
   eoi_flag_reg : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N446, next_state => cmd_26_port, 
               clocked_on => clk_port, Q => eoi_flag, QN => n_1181);
   eot_flag_reg : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N446, next_state => cmd_25_port, 
               clocked_on => clk_port, Q => eot_flag, QN => n_1182);
   keyPISO : KEY_PISO_2 port map( clk => clk_port, rst => rst, data_s(31) => 
                           key(31), data_s(30) => key(30), data_s(29) => 
                           key(29), data_s(28) => key(28), data_s(27) => 
                           key(27), data_s(26) => key(26), data_s(25) => 
                           key(25), data_s(24) => key(24), data_s(23) => 
                           key(23), data_s(22) => key(22), data_s(21) => 
                           key(21), data_s(20) => key(20), data_s(19) => 
                           key(19), data_s(18) => key(18), data_s(17) => 
                           key(17), data_s(16) => key(16), data_s(15) => 
                           key(15), data_s(14) => key(14), data_s(13) => 
                           key(13), data_s(12) => key(12), data_s(11) => 
                           key(11), data_s(10) => key(10), data_s(9) => key(9),
                           data_s(8) => key(8), data_s(7) => key(7), data_s(6) 
                           => key(6), data_s(5) => key(5), data_s(4) => key(4),
                           data_s(3) => key(3), data_s(2) => key(2), data_s(1) 
                           => key(1), data_s(0) => key(0), data_valid_s => 
                           key_valid, data_ready_s => key_ready, data_p(31) => 
                           sdi_data_31_port, data_p(30) => sdi_data_30_port, 
                           data_p(29) => sdi_data_29_port, data_p(28) => 
                           sdi_data_28_port, data_p(27) => sdi_data_27_port, 
                           data_p(26) => sdi_data_26_port, data_p(25) => 
                           sdi_data_25_port, data_p(24) => sdi_data_24_port, 
                           data_p(23) => sdi_data_23_port, data_p(22) => 
                           sdi_data_22_port, data_p(21) => sdi_data_21_port, 
                           data_p(20) => sdi_data_20_port, data_p(19) => 
                           sdi_data_19_port, data_p(18) => sdi_data_18_port, 
                           data_p(17) => sdi_data_17_port, data_p(16) => 
                           sdi_data_16_port, data_p(15) => sdi_data_15_port, 
                           data_p(14) => sdi_data_14_port, data_p(13) => 
                           sdi_data_13_port, data_p(12) => sdi_data_12_port, 
                           data_p(11) => sdi_data_11_port, data_p(10) => 
                           sdi_data_10_port, data_p(9) => sdi_data_9_port, 
                           data_p(8) => sdi_data_8_port, data_p(7) => 
                           sdi_data_7_port, data_p(6) => sdi_data_6_port, 
                           data_p(5) => sdi_data_5_port, data_p(4) => 
                           sdi_data_4_port, data_p(3) => sdi_data_3_port, 
                           data_p(2) => sdi_data_2_port, data_p(1) => 
                           sdi_data_1_port, data_p(0) => sdi_data_0_port, 
                           data_valid_p => key_valid_p, data_ready_p => 
                           key_ready_p);
   bdiPISO : DATA_PISO_2 port map( clk => clk_port, rst => rst, data_size_p(2) 
                           => bdi_size_p_2_port, data_size_p(1) => 
                           bdi_size_p_1_port, data_size_p(0) => 
                           bdi_size_p_0_port, data_size_s(2) => bdi_size(2), 
                           data_size_s(1) => bdi_size(1), data_size_s(0) => 
                           bdi_size(0), data_s(31) => bdi(31), data_s(30) => 
                           bdi(30), data_s(29) => bdi(29), data_s(28) => 
                           bdi(28), data_s(27) => bdi(27), data_s(26) => 
                           bdi(26), data_s(25) => bdi(25), data_s(24) => 
                           bdi(24), data_s(23) => bdi(23), data_s(22) => 
                           bdi(22), data_s(21) => bdi(21), data_s(20) => 
                           bdi(20), data_s(19) => bdi(19), data_s(18) => 
                           bdi(18), data_s(17) => bdi(17), data_s(16) => 
                           bdi(16), data_s(15) => bdi(15), data_s(14) => 
                           bdi(14), data_s(13) => bdi(13), data_s(12) => 
                           bdi(12), data_s(11) => bdi(11), data_s(10) => 
                           bdi(10), data_s(9) => bdi(9), data_s(8) => bdi(8), 
                           data_s(7) => bdi(7), data_s(6) => bdi(6), data_s(5) 
                           => bdi(5), data_s(4) => bdi(4), data_s(3) => bdi(3),
                           data_s(2) => bdi(2), data_s(1) => bdi(1), data_s(0) 
                           => bdi(0), data_valid_s => bdi_valid, data_ready_s 
                           => bdi_ready, data_p(31) => cmd_31_port, data_p(30) 
                           => cmd_30_port, data_p(29) => cmd_29_port, 
                           data_p(28) => cmd_28_port, data_p(27) => cmd_27_port
                           , data_p(26) => cmd_26_port, data_p(25) => 
                           cmd_25_port, data_p(24) => cmd_24_port, data_p(23) 
                           => cmd_23_port, data_p(22) => cmd_22_port, 
                           data_p(21) => cmd_21_port, data_p(20) => cmd_20_port
                           , data_p(19) => cmd_19_port, data_p(18) => 
                           cmd_18_port, data_p(17) => cmd_17_port, data_p(16) 
                           => cmd_16_port, data_p(15) => cmd_15_port, 
                           data_p(14) => cmd_14_port, data_p(13) => cmd_13_port
                           , data_p(12) => cmd_12_port, data_p(11) => 
                           cmd_11_port, data_p(10) => cmd_10_port, data_p(9) =>
                           cmd_9_port, data_p(8) => cmd_8_port, data_p(7) => 
                           cmd_7_port, data_p(6) => cmd_6_port, data_p(5) => 
                           cmd_5_port, data_p(4) => cmd_4_port, data_p(3) => 
                           cmd_3_port, data_p(2) => cmd_2_port, data_p(1) => 
                           cmd_1_port, data_p(0) => cmd_0_port, data_valid_p =>
                           bdi_valid_p, data_ready_p => bdi_ready_p, 
                           valid_bytes_p(3) => bdi_valid_bytes_p_3_port, 
                           valid_bytes_p(2) => bdi_valid_bytes_p_2_port, 
                           valid_bytes_p(1) => bdi_valid_bytes_p_1_port, 
                           valid_bytes_p(0) => bdi_valid_bytes_p_0_port, 
                           valid_bytes_s(3) => bdi_valid_bytes(3), 
                           valid_bytes_s(2) => bdi_valid_bytes(2), 
                           valid_bytes_s(1) => bdi_valid_bytes(1), 
                           valid_bytes_s(0) => bdi_valid_bytes(0), pad_loc_p(3)
                           => bdi_pad_loc_p_3_port, pad_loc_p(2) => 
                           bdi_pad_loc_p_2_port, pad_loc_p(1) => 
                           bdi_pad_loc_p_1_port, pad_loc_p(0) => 
                           bdi_pad_loc_p_0_port, pad_loc_s(3) => bdi_pad_loc(3)
                           , pad_loc_s(2) => bdi_pad_loc(2), pad_loc_s(1) => 
                           bdi_pad_loc(1), pad_loc_s(0) => bdi_pad_loc(0), 
                           eoi_p => bdi_eoi_internal, eoi_s => bdi_eoi, eot_p 
                           => bdi_eot_internal, eot_s => bdi_eot);
   pr_state_reg_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => X_Logic1_port, next_state => N209
               , clocked_on => clk_port, Q => pr_state_3_port, QN => n_1183);
   pr_state_reg_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => X_Logic1_port, next_state => N208
               , clocked_on => clk_port, Q => pr_state_2_port, QN => n_1184);
   pr_state_reg_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => X_Logic1_port, next_state => N207
               , clocked_on => clk_port, Q => pr_state_1_port, QN => n_1185);
   pr_state_reg_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => X_Logic1_port, next_state => N206
               , clocked_on => clk_port, Q => pr_state_0_port, QN => n_1186);
   C230 : GTECH_AND2 port map( A => N210, B => N211, Z => N214);
   C231 : GTECH_AND2 port map( A => N212, B => N213, Z => N215);
   C232 : GTECH_AND2 port map( A => N214, B => N215, Z => N216);
   C234 : GTECH_OR2 port map( A => pr_state_3_port, B => pr_state_2_port, Z => 
                           N217);
   C235 : GTECH_OR2 port map( A => pr_state_1_port, B => N213, Z => N218);
   C236 : GTECH_OR2 port map( A => N217, B => N218, Z => N219);
   C239 : GTECH_OR2 port map( A => pr_state_3_port, B => pr_state_2_port, Z => 
                           N221);
   C240 : GTECH_OR2 port map( A => N212, B => pr_state_0_port, Z => N222);
   C241 : GTECH_OR2 port map( A => N221, B => N222, Z => N223);
   C245 : GTECH_OR2 port map( A => pr_state_3_port, B => pr_state_2_port, Z => 
                           N225);
   C246 : GTECH_OR2 port map( A => N212, B => N213, Z => N226);
   C247 : GTECH_OR2 port map( A => N225, B => N226, Z => N227);
   C250 : GTECH_OR2 port map( A => pr_state_3_port, B => N211, Z => N229);
   C251 : GTECH_OR2 port map( A => pr_state_1_port, B => pr_state_0_port, Z => 
                           N230);
   C252 : GTECH_OR2 port map( A => N229, B => N230, Z => N231);
   C256 : GTECH_OR2 port map( A => pr_state_3_port, B => N211, Z => N233);
   C257 : GTECH_OR2 port map( A => pr_state_1_port, B => N213, Z => N234);
   C258 : GTECH_OR2 port map( A => N233, B => N234, Z => N235);
   C262 : GTECH_OR2 port map( A => pr_state_3_port, B => N211, Z => N237);
   C263 : GTECH_OR2 port map( A => N212, B => pr_state_0_port, Z => N238);
   C264 : GTECH_OR2 port map( A => N237, B => N238, Z => N239);
   C269 : GTECH_OR2 port map( A => pr_state_3_port, B => N211, Z => N241);
   C270 : GTECH_OR2 port map( A => N212, B => N213, Z => N242);
   C271 : GTECH_OR2 port map( A => N241, B => N242, Z => N243);
   C274 : GTECH_OR2 port map( A => N210, B => pr_state_2_port, Z => N245);
   C275 : GTECH_OR2 port map( A => pr_state_1_port, B => pr_state_0_port, Z => 
                           N246);
   C276 : GTECH_OR2 port map( A => N245, B => N246, Z => N247);
   C280 : GTECH_OR2 port map( A => N210, B => pr_state_2_port, Z => N249);
   C281 : GTECH_OR2 port map( A => pr_state_1_port, B => N213, Z => N250);
   C282 : GTECH_OR2 port map( A => N249, B => N250, Z => N251);
   C286 : GTECH_OR2 port map( A => N210, B => pr_state_2_port, Z => N253);
   C287 : GTECH_OR2 port map( A => N212, B => pr_state_0_port, Z => N254);
   C288 : GTECH_OR2 port map( A => N253, B => N254, Z => N255);
   C293 : GTECH_OR2 port map( A => N210, B => pr_state_2_port, Z => N257);
   C294 : GTECH_OR2 port map( A => N212, B => N213, Z => N258);
   C295 : GTECH_OR2 port map( A => N257, B => N258, Z => N259);
   C299 : GTECH_OR2 port map( A => N210, B => N211, Z => N261);
   C300 : GTECH_OR2 port map( A => pr_state_1_port, B => pr_state_0_port, Z => 
                           N262);
   C301 : GTECH_OR2 port map( A => N261, B => N262, Z => N263);
   C306 : GTECH_OR2 port map( A => N210, B => N211, Z => N265);
   C307 : GTECH_OR2 port map( A => pr_state_1_port, B => N213, Z => N266);
   C308 : GTECH_OR2 port map( A => N265, B => N266, Z => N267);
   C313 : GTECH_OR2 port map( A => N210, B => N211, Z => N269);
   C314 : GTECH_OR2 port map( A => N212, B => pr_state_0_port, Z => N270);
   C315 : GTECH_OR2 port map( A => N269, B => N270, Z => N271);
   C317 : GTECH_AND2 port map( A => pr_state_3_port, B => pr_state_2_port, Z =>
                           N273);
   C318 : GTECH_AND2 port map( A => pr_state_1_port, B => pr_state_0_port, Z =>
                           N274);
   C319 : GTECH_AND2 port map( A => N273, B => N274, Z => N275);
   C619 : GTECH_AND2 port map( A => N210, B => N211, Z => N329);
   C620 : GTECH_AND2 port map( A => N212, B => N213, Z => N330);
   C621 : GTECH_AND2 port map( A => N329, B => N330, Z => N331);
   C623 : GTECH_OR2 port map( A => pr_state_3_port, B => pr_state_2_port, Z => 
                           N332);
   C624 : GTECH_OR2 port map( A => pr_state_1_port, B => N213, Z => N333);
   C625 : GTECH_OR2 port map( A => N332, B => N333, Z => N334);
   C628 : GTECH_OR2 port map( A => pr_state_3_port, B => pr_state_2_port, Z => 
                           N336);
   C629 : GTECH_OR2 port map( A => N212, B => pr_state_0_port, Z => N337);
   C630 : GTECH_OR2 port map( A => N336, B => N337, Z => N338);
   C634 : GTECH_OR2 port map( A => pr_state_3_port, B => pr_state_2_port, Z => 
                           N340);
   C635 : GTECH_OR2 port map( A => N212, B => N213, Z => N341);
   C636 : GTECH_OR2 port map( A => N340, B => N341, Z => N342);
   C639 : GTECH_OR2 port map( A => pr_state_3_port, B => N211, Z => N344);
   C640 : GTECH_OR2 port map( A => pr_state_1_port, B => pr_state_0_port, Z => 
                           N345);
   C641 : GTECH_OR2 port map( A => N344, B => N345, Z => N346);
   C645 : GTECH_OR2 port map( A => pr_state_3_port, B => N211, Z => N348);
   C646 : GTECH_OR2 port map( A => pr_state_1_port, B => N213, Z => N349);
   C647 : GTECH_OR2 port map( A => N348, B => N349, Z => N350);
   C651 : GTECH_OR2 port map( A => pr_state_3_port, B => N211, Z => N352);
   C652 : GTECH_OR2 port map( A => N212, B => pr_state_0_port, Z => N353);
   C653 : GTECH_OR2 port map( A => N352, B => N353, Z => N354);
   C658 : GTECH_OR2 port map( A => pr_state_3_port, B => N211, Z => N356);
   C659 : GTECH_OR2 port map( A => N212, B => N213, Z => N357);
   C660 : GTECH_OR2 port map( A => N356, B => N357, Z => N358);
   C663 : GTECH_OR2 port map( A => N210, B => pr_state_2_port, Z => N360);
   C664 : GTECH_OR2 port map( A => pr_state_1_port, B => pr_state_0_port, Z => 
                           N361);
   C665 : GTECH_OR2 port map( A => N360, B => N361, Z => N362);
   C669 : GTECH_OR2 port map( A => N210, B => pr_state_2_port, Z => N364);
   C670 : GTECH_OR2 port map( A => pr_state_1_port, B => N213, Z => N365);
   C671 : GTECH_OR2 port map( A => N364, B => N365, Z => N366);
   C675 : GTECH_OR2 port map( A => N210, B => pr_state_2_port, Z => N368);
   C676 : GTECH_OR2 port map( A => N212, B => pr_state_0_port, Z => N369);
   C677 : GTECH_OR2 port map( A => N368, B => N369, Z => N370);
   C682 : GTECH_OR2 port map( A => N210, B => pr_state_2_port, Z => N372);
   C683 : GTECH_OR2 port map( A => N212, B => N213, Z => N373);
   C684 : GTECH_OR2 port map( A => N372, B => N373, Z => N374);
   C688 : GTECH_OR2 port map( A => N210, B => N211, Z => N376);
   C689 : GTECH_OR2 port map( A => pr_state_1_port, B => pr_state_0_port, Z => 
                           N377);
   C690 : GTECH_OR2 port map( A => N376, B => N377, Z => N378);
   C695 : GTECH_OR2 port map( A => N210, B => N211, Z => N380);
   C696 : GTECH_OR2 port map( A => pr_state_1_port, B => N213, Z => N381);
   C697 : GTECH_OR2 port map( A => N380, B => N381, Z => N382);
   C702 : GTECH_OR2 port map( A => N210, B => N211, Z => N384);
   C703 : GTECH_OR2 port map( A => N212, B => pr_state_0_port, Z => N385);
   C704 : GTECH_OR2 port map( A => N384, B => N385, Z => N386);
   C706 : GTECH_AND2 port map( A => pr_state_3_port, B => pr_state_2_port, Z =>
                           N388);
   C707 : GTECH_AND2 port map( A => pr_state_1_port, B => pr_state_0_port, Z =>
                           N389);
   C708 : GTECH_AND2 port map( A => N388, B => N389, Z => N390);
   I_10 : GTECH_NOT port map( A => cmd_31_port, Z => N447);
   C923 : GTECH_OR2 port map( A => cmd_30_port, B => N447, Z => N448);
   C924 : GTECH_OR2 port map( A => cmd_29_port, B => N448, Z => N449);
   C925 : GTECH_OR2 port map( A => cmd_28_port, B => N449, Z => N450);
   I_11 : GTECH_NOT port map( A => N450, Z => N451);
   C927 : GTECH_OR2 port map( A => cmd_14_port, B => cmd_15_port, Z => N452);
   C928 : GTECH_OR2 port map( A => cmd_13_port, B => N452, Z => N453);
   C929 : GTECH_OR2 port map( A => cmd_12_port, B => N453, Z => N454);
   C930 : GTECH_OR2 port map( A => cmd_11_port, B => N454, Z => N455);
   C931 : GTECH_OR2 port map( A => cmd_10_port, B => N455, Z => N456);
   C932 : GTECH_OR2 port map( A => cmd_9_port, B => N456, Z => N457);
   C933 : GTECH_OR2 port map( A => cmd_8_port, B => N457, Z => N458);
   C934 : GTECH_OR2 port map( A => cmd_7_port, B => N458, Z => N459);
   C935 : GTECH_OR2 port map( A => cmd_6_port, B => N459, Z => N460);
   C936 : GTECH_OR2 port map( A => cmd_5_port, B => N460, Z => N461);
   C937 : GTECH_OR2 port map( A => cmd_4_port, B => N461, Z => N462);
   C938 : GTECH_OR2 port map( A => cmd_3_port, B => N462, Z => N463);
   C939 : GTECH_OR2 port map( A => cmd_2_port, B => N463, Z => N464);
   C940 : GTECH_OR2 port map( A => cmd_1_port, B => N464, Z => N465);
   C941 : GTECH_OR2 port map( A => cmd_0_port, B => N465, Z => N466);
   I_12 : GTECH_NOT port map( A => N466, Z => N467);
   C943 : GTECH_OR2 port map( A => cmd_14_port, B => cmd_15_port, Z => N468);
   C944 : GTECH_OR2 port map( A => cmd_13_port, B => N468, Z => N469);
   C945 : GTECH_OR2 port map( A => cmd_12_port, B => N469, Z => N470);
   C946 : GTECH_OR2 port map( A => cmd_11_port, B => N470, Z => N471);
   C947 : GTECH_OR2 port map( A => cmd_10_port, B => N471, Z => N472);
   C948 : GTECH_OR2 port map( A => cmd_9_port, B => N472, Z => N473);
   C949 : GTECH_OR2 port map( A => cmd_8_port, B => N473, Z => N474);
   C950 : GTECH_OR2 port map( A => cmd_7_port, B => N474, Z => N475);
   C951 : GTECH_OR2 port map( A => cmd_6_port, B => N475, Z => N476);
   C952 : GTECH_OR2 port map( A => cmd_5_port, B => N476, Z => N477);
   C953 : GTECH_OR2 port map( A => cmd_4_port, B => N477, Z => N478);
   C954 : GTECH_OR2 port map( A => cmd_3_port, B => N478, Z => N479);
   C955 : GTECH_OR2 port map( A => cmd_2_port, B => N479, Z => N480);
   C956 : GTECH_OR2 port map( A => cmd_1_port, B => N480, Z => N481);
   C957 : GTECH_OR2 port map( A => cmd_0_port, B => N481, Z => N482);
   I_13 : GTECH_NOT port map( A => N482, Z => N483);
   C959 : GTECH_OR2 port map( A => cmd_14_port, B => cmd_15_port, Z => N484);
   C960 : GTECH_OR2 port map( A => cmd_13_port, B => N484, Z => N485);
   C961 : GTECH_OR2 port map( A => cmd_12_port, B => N485, Z => N486);
   C962 : GTECH_OR2 port map( A => cmd_11_port, B => N486, Z => N487);
   C963 : GTECH_OR2 port map( A => cmd_10_port, B => N487, Z => N488);
   C964 : GTECH_OR2 port map( A => cmd_9_port, B => N488, Z => N489);
   C965 : GTECH_OR2 port map( A => cmd_8_port, B => N489, Z => N490);
   C966 : GTECH_OR2 port map( A => cmd_7_port, B => N490, Z => N491);
   C967 : GTECH_OR2 port map( A => cmd_6_port, B => N491, Z => N492);
   C968 : GTECH_OR2 port map( A => cmd_5_port, B => N492, Z => N493);
   C969 : GTECH_OR2 port map( A => cmd_4_port, B => N493, Z => N494);
   C970 : GTECH_OR2 port map( A => cmd_3_port, B => N494, Z => N495);
   C971 : GTECH_OR2 port map( A => cmd_2_port, B => N495, Z => N496);
   C972 : GTECH_OR2 port map( A => cmd_1_port, B => N496, Z => N497);
   C973 : GTECH_OR2 port map( A => cmd_0_port, B => N497, Z => N498);
   I_14 : GTECH_NOT port map( A => N498, Z => N499);
   C976 : GTECH_OR2 port map( A => cmd_30_port, B => N447, Z => N500);
   C977 : GTECH_OR2 port map( A => cmd_29_port, B => N500, Z => N501);
   C978 : GTECH_OR2 port map( A => cmd_28_port, B => N501, Z => N502);
   I_15 : GTECH_NOT port map( A => N502, Z => N503);
   I_16 : GTECH_NOT port map( A => cmd_29_port, Z => N504);
   C981 : GTECH_OR2 port map( A => cmd_30_port, B => cmd_31_port, Z => N505);
   C982 : GTECH_OR2 port map( A => N504, B => N505, Z => N506);
   C983 : GTECH_OR2 port map( A => cmd_28_port, B => N506, Z => N507);
   I_17 : GTECH_NOT port map( A => N507, Z => N508);
   I_18 : GTECH_NOT port map( A => cmd_28_port, Z => N509);
   C987 : GTECH_OR2 port map( A => cmd_30_port, B => cmd_31_port, Z => N510);
   C988 : GTECH_OR2 port map( A => N504, B => N510, Z => N511);
   C989 : GTECH_OR2 port map( A => N509, B => N511, Z => N512);
   I_19 : GTECH_NOT port map( A => N512, Z => N513);
   C992 : GTECH_OR2 port map( A => cmd_30_port, B => cmd_31_port, Z => N514);
   C993 : GTECH_OR2 port map( A => N504, B => N514, Z => N515);
   C994 : GTECH_OR2 port map( A => cmd_28_port, B => N515, Z => N516);
   I_20 : GTECH_NOT port map( A => N516, Z => N517);
   C998 : GTECH_OR2 port map( A => cmd_30_port, B => cmd_31_port, Z => N518);
   C999 : GTECH_OR2 port map( A => N504, B => N518, Z => N519);
   C1000 : GTECH_OR2 port map( A => N509, B => N519, Z => N520);
   I_21 : GTECH_NOT port map( A => N520, Z => N521);
   I_22 : GTECH_NOT port map( A => cmd_30_port, Z => N522);
   C1005 : GTECH_OR2 port map( A => N522, B => cmd_31_port, Z => N523);
   C1006 : GTECH_OR2 port map( A => N504, B => N523, Z => N524);
   C1007 : GTECH_OR2 port map( A => N509, B => N524, Z => N525);
   I_23 : GTECH_NOT port map( A => N525, Z => N526);
   C1009_cell : SELECT_OP
      generic map ( num_inputs => 5, input_width => 4 )
      port map(
         -- Connections to port 'DATA1'
         DATA(3) => X_Logic0_port, DATA(2) => X_Logic0_port, DATA(1) => 
               X_Logic0_port, DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(7) => X_Logic1_port, DATA(6) => X_Logic0_port, DATA(5) => 
               X_Logic0_port, DATA(4) => X_Logic0_port, 
         -- Connections to port 'DATA3'
         DATA(11) => X_Logic1_port, DATA(10) => X_Logic1_port, DATA(9) => 
               X_Logic0_port, DATA(8) => X_Logic0_port, 
         -- Connections to port 'DATA4'
         DATA(15) => X_Logic1_port, DATA(14) => X_Logic1_port, DATA(13) => 
               X_Logic1_port, DATA(12) => X_Logic0_port, 
         -- Connections to port 'DATA5'
         DATA(19) => X_Logic1_port, DATA(18) => X_Logic1_port, DATA(17) => 
               X_Logic1_port, DATA(16) => X_Logic1_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N0, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N1, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N2, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N3, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N134, 
         -- Connections to port 'Z'
         Z(3) => bdi_valid_bytes_p_3_port, Z(2) => bdi_valid_bytes_p_2_port, 
               Z(1) => bdi_valid_bytes_p_1_port, Z(0) => 
               bdi_valid_bytes_p_0_port );
   B_0 : GTECH_BUF port map( A => N80, Z => N0);
   B_1 : GTECH_BUF port map( A => N97, Z => N1);
   B_2 : GTECH_BUF port map( A => N114, Z => N2);
   B_3 : GTECH_BUF port map( A => N130, Z => N3);
   C1010_cell : SELECT_OP
      generic map ( num_inputs => 5, input_width => 4 )
      port map(
         -- Connections to port 'DATA1'
         DATA(3) => X_Logic1_port, DATA(2) => X_Logic0_port, DATA(1) => 
               X_Logic0_port, DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(7) => X_Logic0_port, DATA(6) => X_Logic1_port, DATA(5) => 
               X_Logic0_port, DATA(4) => X_Logic0_port, 
         -- Connections to port 'DATA3'
         DATA(11) => X_Logic0_port, DATA(10) => X_Logic0_port, DATA(9) => 
               X_Logic1_port, DATA(8) => X_Logic0_port, 
         -- Connections to port 'DATA4'
         DATA(15) => X_Logic0_port, DATA(14) => X_Logic0_port, DATA(13) => 
               X_Logic0_port, DATA(12) => X_Logic1_port, 
         -- Connections to port 'DATA5'
         DATA(19) => X_Logic0_port, DATA(18) => X_Logic0_port, DATA(17) => 
               X_Logic0_port, DATA(16) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N4, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N5, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N6, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N7, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N202, 
         -- Connections to port 'Z'
         Z(3) => bdi_pad_loc_p_3_port, Z(2) => bdi_pad_loc_p_2_port, Z(1) => 
               bdi_pad_loc_p_1_port, Z(0) => bdi_pad_loc_p_0_port );
   B_4 : GTECH_BUF port map( A => N150, Z => N4);
   B_5 : GTECH_BUF port map( A => N166, Z => N5);
   B_6 : GTECH_BUF port map( A => N182, Z => N6);
   B_7 : GTECH_BUF port map( A => N198, Z => N7);
   C1011_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 16 )
      port map(
         -- Connections to port 'DATA1'
         DATA(15) => sdi_data_15_port, DATA(14) => sdi_data_14_port, DATA(13) 
               => sdi_data_13_port, DATA(12) => sdi_data_12_port, DATA(11) => 
               sdi_data_11_port, DATA(10) => sdi_data_10_port, DATA(9) => 
               sdi_data_9_port, DATA(8) => sdi_data_8_port, DATA(7) => 
               sdi_data_7_port, DATA(6) => sdi_data_6_port, DATA(5) => 
               sdi_data_5_port, DATA(4) => sdi_data_4_port, DATA(3) => 
               sdi_data_3_port, DATA(2) => sdi_data_2_port, DATA(1) => 
               sdi_data_1_port, DATA(0) => sdi_data_0_port, 
         -- Connections to port 'DATA2'
         DATA(31) => cmd_15_port, DATA(30) => cmd_14_port, DATA(29) => 
               cmd_13_port, DATA(28) => cmd_12_port, DATA(27) => cmd_11_port, 
               DATA(26) => cmd_10_port, DATA(25) => cmd_9_port, DATA(24) => 
               cmd_8_port, DATA(23) => cmd_7_port, DATA(22) => cmd_6_port, 
               DATA(21) => cmd_5_port, DATA(20) => cmd_4_port, DATA(19) => 
               cmd_3_port, DATA(18) => cmd_2_port, DATA(17) => cmd_1_port, 
               DATA(16) => cmd_0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N8, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N9, 
         -- Connections to port 'Z'
         Z(15) => load_SegLenCnt_15_port, Z(14) => load_SegLenCnt_14_port, 
               Z(13) => load_SegLenCnt_13_port, Z(12) => load_SegLenCnt_12_port
               , Z(11) => load_SegLenCnt_11_port, Z(10) => 
               load_SegLenCnt_10_port, Z(9) => load_SegLenCnt_9_port, Z(8) => 
               load_SegLenCnt_8_port, Z(7) => load_SegLenCnt_7_port, Z(6) => 
               load_SegLenCnt_6_port, Z(5) => load_SegLenCnt_5_port, Z(4) => 
               load_SegLenCnt_4_port, Z(3) => load_SegLenCnt_3_port, Z(2) => 
               load_SegLenCnt_2_port, Z(1) => load_SegLenCnt_1_port, Z(0) => 
               load_SegLenCnt_0_port );
   B_8 : GTECH_BUF port map( A => sel_sdi_length, Z => N8);
   B_9 : GTECH_BUF port map( A => N203, Z => N9);
   C1012_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 3 )
      port map(
         -- Connections to port 'DATA1'
         DATA(2) => dout_SegLenCnt_2_port, DATA(1) => dout_SegLenCnt_1_port, 
               DATA(0) => dout_SegLenCnt_0_port, 
         -- Connections to port 'DATA2'
         DATA(5) => X_Logic1_port, DATA(4) => X_Logic0_port, DATA(3) => 
               X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N10, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N11, 
         -- Connections to port 'Z'
         Z(2) => bdi_size_p_2_port, Z(1) => bdi_size_p_1_port, Z(0) => 
               bdi_size_p_0_port );
   B_10 : GTECH_BUF port map( A => last_flit_of_segment, Z => N10);
   B_11 : GTECH_BUF port map( A => N204, Z => N11);
   C1013_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 4 )
      port map(
         -- Connections to port 'DATA1'
         DATA(3) => X_Logic0_port, DATA(2) => X_Logic0_port, DATA(1) => 
               X_Logic0_port, DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(7) => nx_state_3_port, DATA(6) => nx_state_2_port, DATA(5) => 
               nx_state_1_port, DATA(4) => nx_state_0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N12, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N13, 
         -- Connections to port 'Z'
         Z(3) => N209, Z(2) => N208, Z(1) => N207, Z(0) => N206 );
   B_12 : GTECH_BUF port map( A => rst, Z => N12);
   B_13 : GTECH_BUF port map( A => N205, Z => N13);
   C1014_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 2 )
      port map(
         -- Connections to port 'DATA1'
         DATA(1) => X_Logic0_port, DATA(0) => X_Logic1_port, 
         -- Connections to port 'DATA2'
         DATA(3) => N278, DATA(2) => N278, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N14, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N277, 
         -- Connections to port 'Z'
         Z(1) => N280, Z(0) => N279 );
   B_14 : GTECH_BUF port map( A => N276, Z => N14);
   C1015_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 2 )
      port map(
         -- Connections to port 'DATA1'
         DATA(1) => X_Logic0_port, DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(3) => N280, DATA(2) => N279, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N15, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N16, 
         -- Connections to port 'Z'
         Z(1) => N282, Z(0) => N281 );
   B_15 : GTECH_BUF port map( A => N526, Z => N15);
   B_16 : GTECH_BUF port map( A => N525, Z => N16);
   C1016_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 3 )
      port map(
         -- Connections to port 'DATA1'
         DATA(2) => N282, DATA(1) => N281, DATA(0) => N526, 
         -- Connections to port 'DATA2'
         DATA(5) => X_Logic0_port, DATA(4) => X_Logic0_port, DATA(3) => 
               X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N17, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N18, 
         -- Connections to port 'Z'
         Z(2) => N285, Z(1) => N284, Z(0) => N283 );
   B_17 : GTECH_BUF port map( A => pdi_valid_port, Z => N17);
   B_18 : GTECH_BUF port map( A => N393, Z => N18);
   I_24 : GTECH_NOT port map( A => N287, Z => N288);
   I_25 : GTECH_NOT port map( A => N289, Z => N290);
   I_26 : GTECH_NOT port map( A => N291, Z => N292);
   C1020_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 3 )
      port map(
         -- Connections to port 'DATA1'
         DATA(2) => N291, DATA(1) => N292, DATA(0) => N292, 
         -- Connections to port 'DATA2'
         DATA(5) => X_Logic0_port, DATA(4) => X_Logic1_port, DATA(3) => 
               X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N17, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N18, 
         -- Connections to port 'Z'
         Z(2) => N295, Z(1) => N294, Z(0) => N293 );
   I_27 : GTECH_NOT port map( A => N296, Z => N299);
   C1022_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 2 )
      port map(
         -- Connections to port 'DATA1'
         DATA(1) => eot_flag, DATA(0) => N298, 
         -- Connections to port 'DATA2'
         DATA(3) => X_Logic0_port, DATA(2) => X_Logic1_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N19, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N297, 
         -- Connections to port 'Z'
         Z(1) => N301, Z(0) => N300 );
   B_19 : GTECH_BUF port map( A => N296, Z => N19);
   I_28 : GTECH_NOT port map( A => N304, Z => N306);
   C1024_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 2 )
      port map(
         -- Connections to port 'DATA1'
         DATA(1) => decrypt_port, DATA(0) => decrypt_port, 
         -- Connections to port 'DATA2'
         DATA(3) => X_Logic1_port, DATA(2) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N20, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N305, 
         -- Connections to port 'Z'
         Z(1) => N308, Z(0) => N307 );
   B_20 : GTECH_BUF port map( A => N304, Z => N20);
   C1025_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 3 )
      port map(
         -- Connections to port 'DATA1'
         DATA(2) => N308, DATA(1) => N307, DATA(0) => N306, 
         -- Connections to port 'DATA2'
         DATA(5) => X_Logic1_port, DATA(4) => X_Logic0_port, DATA(3) => 
               X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N21, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N303, 
         -- Connections to port 'Z'
         Z(2) => N311, Z(1) => N310, Z(0) => N309 );
   B_21 : GTECH_BUF port map( A => N302, Z => N21);
   C1026_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 2 )
      port map(
         -- Connections to port 'DATA1'
         DATA(1) => decrypt_port, DATA(0) => decrypt_port, 
         -- Connections to port 'DATA2'
         DATA(3) => X_Logic1_port, DATA(2) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N22, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N23, 
         -- Connections to port 'Z'
         Z(1) => N315, Z(0) => N314 );
   B_22 : GTECH_BUF port map( A => eot_flag, Z => N22);
   B_23 : GTECH_BUF port map( A => N298, Z => N23);
   I_29 : GTECH_NOT port map( A => N312, Z => N316);
   C1028_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 2 )
      port map(
         -- Connections to port 'DATA1'
         DATA(1) => N315, DATA(0) => N314, 
         -- Connections to port 'DATA2'
         DATA(3) => X_Logic1_port, DATA(2) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N24, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N313, 
         -- Connections to port 'Z'
         Z(1) => N318, Z(0) => N317 );
   B_24 : GTECH_BUF port map( A => N312, Z => N24);
   C1029_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => N328, 
         -- Connections to port 'DATA2'
         DATA(1) => X_Logic1_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N25, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N320, 
         -- Connections to port 'Z'
         Z(0) => N321 );
   B_25 : GTECH_BUF port map( A => N319, Z => N25);
   C1031_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 2 )
      port map(
         -- Connections to port 'DATA1'
         DATA(1) => N467, DATA(0) => N466, 
         -- Connections to port 'DATA2'
         DATA(3) => X_Logic0_port, DATA(2) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N17, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N18, 
         -- Connections to port 'Z'
         Z(1) => N323, Z(0) => N322 );
   I_30 : GTECH_NOT port map( A => N324, Z => N326);
   C1033_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => N298, 
         -- Connections to port 'DATA2'
         DATA(1) => X_Logic1_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N26, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N325, 
         -- Connections to port 'Z'
         Z(0) => N327 );
   B_26 : GTECH_BUF port map( A => N324, Z => N26);
   C1034_cell : SELECT_OP
      generic map ( num_inputs => 16, input_width => 4 )
      port map(
         -- Connections to port 'DATA1'
         DATA(3) => N285, DATA(2) => N284, DATA(1) => X_Logic0_port, DATA(0) =>
               N283, 
         -- Connections to port 'DATA2'
         DATA(7) => X_Logic0_port, DATA(6) => X_Logic0_port, DATA(5) => 
               sdi_valid_port, DATA(4) => N286, 
         -- Connections to port 'DATA3'
         DATA(11) => X_Logic0_port, DATA(10) => X_Logic0_port, DATA(9) => 
               X_Logic1_port, DATA(8) => sdi_valid_port, 
         -- Connections to port 'DATA4'
         DATA(15) => X_Logic0_port, DATA(14) => X_Logic0_port, DATA(13) => N288
               , DATA(12) => N288, 
         -- Connections to port 'DATA5'
         DATA(19) => X_Logic0_port, DATA(18) => X_Logic1_port, DATA(17) => 
               X_Logic0_port, DATA(16) => pdi_valid_port, 
         -- Connections to port 'DATA6'
         DATA(23) => X_Logic0_port, DATA(22) => X_Logic1_port, DATA(21) => N289
               , DATA(20) => N290, 
         -- Connections to port 'DATA7'
         DATA(27) => N295, DATA(26) => N294, DATA(25) => N294, DATA(24) => N293
               , 
         -- Connections to port 'DATA8'
         DATA(31) => N301, DATA(30) => N300, DATA(29) => N300, DATA(28) => N299
               , 
         -- Connections to port 'DATA9'
         DATA(35) => N311, DATA(34) => X_Logic0_port, DATA(33) => N310, 
               DATA(32) => N309, 
         -- Connections to port 'DATA10'
         DATA(39) => N318, DATA(38) => X_Logic0_port, DATA(37) => N317, 
               DATA(36) => N316, 
         -- Connections to port 'DATA11'
         DATA(43) => X_Logic1_port, DATA(42) => X_Logic0_port, DATA(41) => 
               X_Logic1_port, DATA(40) => pdi_valid_port, 
         -- Connections to port 'DATA12'
         DATA(47) => N321, DATA(46) => X_Logic0_port, DATA(45) => N321, 
               DATA(44) => N321, 
         -- Connections to port 'DATA13'
         DATA(51) => X_Logic1_port, DATA(50) => X_Logic1_port, DATA(49) => N323
               , DATA(48) => N322, 
         -- Connections to port 'DATA14'
         DATA(55) => N327, DATA(54) => N327, DATA(53) => X_Logic0_port, 
               DATA(52) => N326, 
         -- Connections to port 'DATA15'
         DATA(59) => N328, DATA(58) => N328, DATA(57) => N328, DATA(56) => 
               X_Logic0_port, 
         -- Connections to port 'DATA16'
         DATA(63) => X_Logic0_port, DATA(62) => X_Logic0_port, DATA(61) => 
               X_Logic0_port, DATA(60) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N27, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N28, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N29, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N30, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N31, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N32, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N33, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N34, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N35, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N36, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N37, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N38, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N39, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N40, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N41, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N42, 
         -- Connections to port 'Z'
         Z(3) => nx_state_3_port, Z(2) => nx_state_2_port, Z(1) => 
               nx_state_1_port, Z(0) => nx_state_0_port );
   B_27 : GTECH_BUF port map( A => N216, Z => N27);
   B_28 : GTECH_BUF port map( A => N220, Z => N28);
   B_29 : GTECH_BUF port map( A => N224, Z => N29);
   B_30 : GTECH_BUF port map( A => N228, Z => N30);
   B_31 : GTECH_BUF port map( A => N232, Z => N31);
   B_32 : GTECH_BUF port map( A => N236, Z => N32);
   B_33 : GTECH_BUF port map( A => N240, Z => N33);
   B_34 : GTECH_BUF port map( A => N244, Z => N34);
   B_35 : GTECH_BUF port map( A => N248, Z => N35);
   B_36 : GTECH_BUF port map( A => N252, Z => N36);
   B_37 : GTECH_BUF port map( A => N256, Z => N37);
   B_38 : GTECH_BUF port map( A => N260, Z => N38);
   B_39 : GTECH_BUF port map( A => N264, Z => N39);
   B_40 : GTECH_BUF port map( A => N268, Z => N40);
   B_41 : GTECH_BUF port map( A => N272, Z => N41);
   B_42 : GTECH_BUF port map( A => N275, Z => N42);
   C1035_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => cmd_28_port, 
         -- Connections to port 'DATA2'
         DATA(1) => decrypt_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N17, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N18, 
         -- Connections to port 'Z'
         Z(0) => N394 );
   C1036_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => cmd_ready_port, 
         -- Connections to port 'DATA2'
         DATA(1) => X_Logic1_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N17, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N18, 
         -- Connections to port 'Z'
         Z(0) => N395 );
   C1037_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => N395, 
         -- Connections to port 'DATA2'
         DATA(1) => X_Logic1_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N43, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N44, 
         -- Connections to port 'Z'
         Z(0) => N396 );
   B_43 : GTECH_BUF port map( A => N451, Z => N43);
   B_44 : GTECH_BUF port map( A => N450, Z => N44);
   C1038_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => pdi_valid_port, 
         -- Connections to port 'DATA2'
         DATA(1) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N43, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N44, 
         -- Connections to port 'Z'
         Z(0) => N397 );
   C1039_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => N395, 
         -- Connections to port 'DATA2'
         DATA(1) => N396, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N45, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N392, 
         -- Connections to port 'Z'
         Z(0) => N398 );
   B_45 : GTECH_BUF port map( A => N391, Z => N45);
   C1040_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => N394, 
         -- Connections to port 'DATA2'
         DATA(1) => decrypt_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N45, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N392, 
         -- Connections to port 'Z'
         Z(0) => N399 );
   C1041_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => pdi_valid_port, 
         -- Connections to port 'DATA2'
         DATA(1) => N397, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N45, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N392, 
         -- Connections to port 'Z'
         Z(0) => N400 );
   C1042_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => N397, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N45, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N392, 
         -- Connections to port 'Z'
         Z(0) => N401 );
   C1043_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => pdi_valid_port, 
         -- Connections to port 'DATA2'
         DATA(1) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N46, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N47, 
         -- Connections to port 'Z'
         Z(0) => N408 );
   B_46 : GTECH_BUF port map( A => decrypt_port, Z => N46);
   B_47 : GTECH_BUF port map( A => N406, Z => N47);
   C1044_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => bdi_ready_p, 
         -- Connections to port 'DATA2'
         DATA(1) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N46, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N47, 
         -- Connections to port 'Z'
         Z(0) => N409 );
   C1045_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => N407, 
         -- Connections to port 'DATA2'
         DATA(1) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N46, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N47, 
         -- Connections to port 'Z'
         Z(0) => N410 );
   C1046_cell : SELECT_OP
      generic map ( num_inputs => 16, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => N398, 
         -- Connections to port 'DATA2'
         DATA(1) => X_Logic0_port, 
         -- Connections to port 'DATA3'
         DATA(2) => X_Logic0_port, 
         -- Connections to port 'DATA4'
         DATA(3) => X_Logic0_port, 
         -- Connections to port 'DATA5'
         DATA(4) => X_Logic1_port, 
         -- Connections to port 'DATA6'
         DATA(5) => bdi_ready_p, 
         -- Connections to port 'DATA7'
         DATA(6) => X_Logic1_port, 
         -- Connections to port 'DATA8'
         DATA(7) => bdi_ready_p, 
         -- Connections to port 'DATA9'
         DATA(8) => cmd_ready_port, 
         -- Connections to port 'DATA10'
         DATA(9) => bdi_ready_p, 
         -- Connections to port 'DATA11'
         DATA(10) => X_Logic1_port, 
         -- Connections to port 'DATA12'
         DATA(11) => N409, 
         -- Connections to port 'DATA13'
         DATA(12) => X_Logic1_port, 
         -- Connections to port 'DATA14'
         DATA(13) => bdi_ready_p, 
         -- Connections to port 'DATA15'
         DATA(14) => X_Logic0_port, 
         -- Connections to port 'DATA16'
         DATA(15) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N48, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N49, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N50, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N51, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N52, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N53, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N54, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N55, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N56, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N57, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N58, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N59, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N60, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N61, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N62, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N63, 
         -- Connections to port 'Z'
         Z(0) => pdi_ready_port );
   B_48 : GTECH_BUF port map( A => N331, Z => N48);
   B_49 : GTECH_BUF port map( A => N335, Z => N49);
   B_50 : GTECH_BUF port map( A => N339, Z => N50);
   B_51 : GTECH_BUF port map( A => N343, Z => N51);
   B_52 : GTECH_BUF port map( A => N347, Z => N52);
   B_53 : GTECH_BUF port map( A => N351, Z => N53);
   B_54 : GTECH_BUF port map( A => N355, Z => N54);
   B_55 : GTECH_BUF port map( A => N359, Z => N55);
   B_56 : GTECH_BUF port map( A => N363, Z => N56);
   B_57 : GTECH_BUF port map( A => N367, Z => N57);
   B_58 : GTECH_BUF port map( A => N371, Z => N58);
   B_59 : GTECH_BUF port map( A => N375, Z => N59);
   B_60 : GTECH_BUF port map( A => N379, Z => N60);
   B_61 : GTECH_BUF port map( A => N383, Z => N61);
   B_62 : GTECH_BUF port map( A => N387, Z => N62);
   B_63 : GTECH_BUF port map( A => N390, Z => N63);
   C1047_cell : SELECT_OP
      generic map ( num_inputs => 16, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => N400, 
         -- Connections to port 'DATA2'
         DATA(1) => X_Logic0_port, 
         -- Connections to port 'DATA3'
         DATA(2) => X_Logic0_port, 
         -- Connections to port 'DATA4'
         DATA(3) => X_Logic0_port, 
         -- Connections to port 'DATA5'
         DATA(4) => X_Logic0_port, 
         -- Connections to port 'DATA6'
         DATA(5) => X_Logic0_port, 
         -- Connections to port 'DATA7'
         DATA(6) => X_Logic0_port, 
         -- Connections to port 'DATA8'
         DATA(7) => X_Logic0_port, 
         -- Connections to port 'DATA9'
         DATA(8) => pdi_valid_port, 
         -- Connections to port 'DATA10'
         DATA(9) => X_Logic0_port, 
         -- Connections to port 'DATA11'
         DATA(10) => X_Logic0_port, 
         -- Connections to port 'DATA12'
         DATA(11) => X_Logic0_port, 
         -- Connections to port 'DATA13'
         DATA(12) => X_Logic0_port, 
         -- Connections to port 'DATA14'
         DATA(13) => X_Logic0_port, 
         -- Connections to port 'DATA15'
         DATA(14) => X_Logic0_port, 
         -- Connections to port 'DATA16'
         DATA(15) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N48, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N49, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N50, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N51, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N52, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N53, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N54, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N55, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N56, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N57, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N58, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N59, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N60, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N61, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N62, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N63, 
         -- Connections to port 'Z'
         Z(0) => cmd_valid_port );
   C1048_cell : SELECT_OP
      generic map ( num_inputs => 16, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => X_Logic1_port, 
         -- Connections to port 'DATA3'
         DATA(2) => X_Logic1_port, 
         -- Connections to port 'DATA4'
         DATA(3) => key_ready_p, 
         -- Connections to port 'DATA5'
         DATA(4) => X_Logic0_port, 
         -- Connections to port 'DATA6'
         DATA(5) => X_Logic0_port, 
         -- Connections to port 'DATA7'
         DATA(6) => X_Logic0_port, 
         -- Connections to port 'DATA8'
         DATA(7) => X_Logic0_port, 
         -- Connections to port 'DATA9'
         DATA(8) => X_Logic0_port, 
         -- Connections to port 'DATA10'
         DATA(9) => X_Logic0_port, 
         -- Connections to port 'DATA11'
         DATA(10) => X_Logic0_port, 
         -- Connections to port 'DATA12'
         DATA(11) => X_Logic0_port, 
         -- Connections to port 'DATA13'
         DATA(12) => X_Logic0_port, 
         -- Connections to port 'DATA14'
         DATA(13) => X_Logic0_port, 
         -- Connections to port 'DATA15'
         DATA(14) => X_Logic0_port, 
         -- Connections to port 'DATA16'
         DATA(15) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N48, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N49, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N50, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N51, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N52, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N53, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N54, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N55, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N56, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N57, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N58, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N59, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N60, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N61, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N62, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N63, 
         -- Connections to port 'Z'
         Z(0) => sdi_ready_port );
   C1049_cell : SELECT_OP
      generic map ( num_inputs => 16, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => X_Logic0_port, 
         -- Connections to port 'DATA3'
         DATA(2) => X_Logic0_port, 
         -- Connections to port 'DATA4'
         DATA(3) => X_Logic1_port, 
         -- Connections to port 'DATA5'
         DATA(4) => X_Logic0_port, 
         -- Connections to port 'DATA6'
         DATA(5) => X_Logic0_port, 
         -- Connections to port 'DATA7'
         DATA(6) => X_Logic0_port, 
         -- Connections to port 'DATA8'
         DATA(7) => X_Logic0_port, 
         -- Connections to port 'DATA9'
         DATA(8) => X_Logic0_port, 
         -- Connections to port 'DATA10'
         DATA(9) => X_Logic0_port, 
         -- Connections to port 'DATA11'
         DATA(10) => X_Logic0_port, 
         -- Connections to port 'DATA12'
         DATA(11) => X_Logic0_port, 
         -- Connections to port 'DATA13'
         DATA(12) => X_Logic0_port, 
         -- Connections to port 'DATA14'
         DATA(13) => X_Logic0_port, 
         -- Connections to port 'DATA15'
         DATA(14) => X_Logic0_port, 
         -- Connections to port 'DATA16'
         DATA(15) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N48, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N49, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N50, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N51, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N52, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N53, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N54, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N55, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N56, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N57, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N58, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N59, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N60, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N61, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N62, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N63, 
         -- Connections to port 'Z'
         Z(0) => key_update_port );
   C1050_cell : SELECT_OP
      generic map ( num_inputs => 16, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => X_Logic0_port, 
         -- Connections to port 'DATA3'
         DATA(2) => sdi_valid_port, 
         -- Connections to port 'DATA4'
         DATA(3) => X_Logic0_port, 
         -- Connections to port 'DATA5'
         DATA(4) => pdi_valid_port, 
         -- Connections to port 'DATA6'
         DATA(5) => X_Logic0_port, 
         -- Connections to port 'DATA7'
         DATA(6) => pdi_valid_port, 
         -- Connections to port 'DATA8'
         DATA(7) => X_Logic0_port, 
         -- Connections to port 'DATA9'
         DATA(8) => N302, 
         -- Connections to port 'DATA10'
         DATA(9) => X_Logic0_port, 
         -- Connections to port 'DATA11'
         DATA(10) => pdi_valid_port, 
         -- Connections to port 'DATA12'
         DATA(11) => X_Logic0_port, 
         -- Connections to port 'DATA13'
         DATA(12) => pdi_valid_port, 
         -- Connections to port 'DATA14'
         DATA(13) => X_Logic0_port, 
         -- Connections to port 'DATA15'
         DATA(14) => X_Logic0_port, 
         -- Connections to port 'DATA16'
         DATA(15) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N48, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N49, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N50, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N51, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N52, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N53, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N54, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N55, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N56, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N57, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N58, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N59, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N60, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N61, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N62, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N63, 
         -- Connections to port 'Z'
         Z(0) => len_SegLenCnt );
   C1051_cell : SELECT_OP
      generic map ( num_inputs => 16, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => X_Logic0_port, 
         -- Connections to port 'DATA3'
         DATA(2) => X_Logic1_port, 
         -- Connections to port 'DATA4'
         DATA(3) => X_Logic0_port, 
         -- Connections to port 'DATA5'
         DATA(4) => X_Logic0_port, 
         -- Connections to port 'DATA6'
         DATA(5) => X_Logic0_port, 
         -- Connections to port 'DATA7'
         DATA(6) => X_Logic0_port, 
         -- Connections to port 'DATA8'
         DATA(7) => X_Logic0_port, 
         -- Connections to port 'DATA9'
         DATA(8) => X_Logic0_port, 
         -- Connections to port 'DATA10'
         DATA(9) => X_Logic0_port, 
         -- Connections to port 'DATA11'
         DATA(10) => X_Logic0_port, 
         -- Connections to port 'DATA12'
         DATA(11) => X_Logic0_port, 
         -- Connections to port 'DATA13'
         DATA(12) => X_Logic0_port, 
         -- Connections to port 'DATA14'
         DATA(13) => X_Logic0_port, 
         -- Connections to port 'DATA15'
         DATA(14) => X_Logic0_port, 
         -- Connections to port 'DATA16'
         DATA(15) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N48, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N49, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N50, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N51, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N52, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N53, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N54, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N55, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N56, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N57, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N58, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N59, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N60, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N61, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N62, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N63, 
         -- Connections to port 'Z'
         Z(0) => sel_sdi_length );
   C1052_cell : SELECT_OP
      generic map ( num_inputs => 16, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => X_Logic0_port, 
         -- Connections to port 'DATA3'
         DATA(2) => X_Logic0_port, 
         -- Connections to port 'DATA4'
         DATA(3) => sdi_valid_port, 
         -- Connections to port 'DATA5'
         DATA(4) => X_Logic0_port, 
         -- Connections to port 'DATA6'
         DATA(5) => X_Logic0_port, 
         -- Connections to port 'DATA7'
         DATA(6) => X_Logic0_port, 
         -- Connections to port 'DATA8'
         DATA(7) => X_Logic0_port, 
         -- Connections to port 'DATA9'
         DATA(8) => X_Logic0_port, 
         -- Connections to port 'DATA10'
         DATA(9) => X_Logic0_port, 
         -- Connections to port 'DATA11'
         DATA(10) => X_Logic0_port, 
         -- Connections to port 'DATA12'
         DATA(11) => X_Logic0_port, 
         -- Connections to port 'DATA13'
         DATA(12) => X_Logic0_port, 
         -- Connections to port 'DATA14'
         DATA(13) => X_Logic0_port, 
         -- Connections to port 'DATA15'
         DATA(14) => X_Logic0_port, 
         -- Connections to port 'DATA16'
         DATA(15) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N48, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N49, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N50, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N51, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N52, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N53, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N54, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N55, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N56, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N57, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N58, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N59, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N60, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N61, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N62, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N63, 
         -- Connections to port 'Z'
         Z(0) => key_valid_p );
   C1053_cell : SELECT_OP
      generic map ( num_inputs => 16, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => X_Logic0_port, 
         -- Connections to port 'DATA3'
         DATA(2) => X_Logic0_port, 
         -- Connections to port 'DATA4'
         DATA(3) => N402, 
         -- Connections to port 'DATA5'
         DATA(4) => X_Logic0_port, 
         -- Connections to port 'DATA6'
         DATA(5) => N403, 
         -- Connections to port 'DATA7'
         DATA(6) => X_Logic0_port, 
         -- Connections to port 'DATA8'
         DATA(7) => N404, 
         -- Connections to port 'DATA9'
         DATA(8) => X_Logic0_port, 
         -- Connections to port 'DATA10'
         DATA(9) => N405, 
         -- Connections to port 'DATA11'
         DATA(10) => X_Logic0_port, 
         -- Connections to port 'DATA12'
         DATA(11) => N410, 
         -- Connections to port 'DATA13'
         DATA(12) => X_Logic0_port, 
         -- Connections to port 'DATA14'
         DATA(13) => N411, 
         -- Connections to port 'DATA15'
         DATA(14) => X_Logic0_port, 
         -- Connections to port 'DATA16'
         DATA(15) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N48, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N49, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N50, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N51, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N52, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N53, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N54, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N55, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N56, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N57, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N58, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N59, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N60, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N61, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N62, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N63, 
         -- Connections to port 'Z'
         Z(0) => en_SegLenCnt );
   C1054_cell : SELECT_OP
      generic map ( num_inputs => 16, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(1) => X_Logic0_port, 
         -- Connections to port 'DATA3'
         DATA(2) => X_Logic0_port, 
         -- Connections to port 'DATA4'
         DATA(3) => X_Logic0_port, 
         -- Connections to port 'DATA5'
         DATA(4) => X_Logic0_port, 
         -- Connections to port 'DATA6'
         DATA(5) => pdi_valid_port, 
         -- Connections to port 'DATA7'
         DATA(6) => X_Logic0_port, 
         -- Connections to port 'DATA8'
         DATA(7) => pdi_valid_port, 
         -- Connections to port 'DATA9'
         DATA(8) => X_Logic0_port, 
         -- Connections to port 'DATA10'
         DATA(9) => pdi_valid_port, 
         -- Connections to port 'DATA11'
         DATA(10) => X_Logic0_port, 
         -- Connections to port 'DATA12'
         DATA(11) => N408, 
         -- Connections to port 'DATA13'
         DATA(12) => X_Logic0_port, 
         -- Connections to port 'DATA14'
         DATA(13) => pdi_valid_port, 
         -- Connections to port 'DATA15'
         DATA(14) => X_Logic1_port, 
         -- Connections to port 'DATA16'
         DATA(15) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N48, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N49, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N50, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N51, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N52, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N53, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N54, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N55, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N56, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N57, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N58, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N59, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N60, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N61, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N62, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N63, 
         -- Connections to port 'Z'
         Z(0) => bdi_valid_p );
   C1055_cell : SELECT_OP
      generic map ( num_inputs => 16, input_width => 4 )
      port map(
         -- Connections to port 'DATA1'
         DATA(3) => X_Logic0_port, DATA(2) => X_Logic0_port, DATA(1) => 
               X_Logic0_port, DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(7) => X_Logic0_port, DATA(6) => X_Logic0_port, DATA(5) => 
               X_Logic0_port, DATA(4) => X_Logic0_port, 
         -- Connections to port 'DATA3'
         DATA(11) => X_Logic0_port, DATA(10) => X_Logic0_port, DATA(9) => 
               X_Logic0_port, DATA(8) => X_Logic0_port, 
         -- Connections to port 'DATA4'
         DATA(15) => X_Logic0_port, DATA(14) => X_Logic0_port, DATA(13) => 
               X_Logic0_port, DATA(12) => X_Logic0_port, 
         -- Connections to port 'DATA5'
         DATA(19) => X_Logic0_port, DATA(18) => X_Logic0_port, DATA(17) => 
               X_Logic0_port, DATA(16) => X_Logic0_port, 
         -- Connections to port 'DATA6'
         DATA(23) => X_Logic1_port, DATA(22) => X_Logic1_port, DATA(21) => 
               X_Logic0_port, DATA(20) => X_Logic1_port, 
         -- Connections to port 'DATA7'
         DATA(27) => X_Logic0_port, DATA(26) => X_Logic0_port, DATA(25) => 
               X_Logic0_port, DATA(24) => X_Logic0_port, 
         -- Connections to port 'DATA8'
         DATA(31) => X_Logic0_port, DATA(30) => X_Logic0_port, DATA(29) => 
               X_Logic0_port, DATA(28) => X_Logic1_port, 
         -- Connections to port 'DATA9'
         DATA(35) => X_Logic0_port, DATA(34) => X_Logic0_port, DATA(33) => 
               X_Logic0_port, DATA(32) => X_Logic0_port, 
         -- Connections to port 'DATA10'
         DATA(39) => X_Logic0_port, DATA(38) => X_Logic1_port, DATA(37) => 
               X_Logic0_port, DATA(36) => decrypt_port, 
         -- Connections to port 'DATA11'
         DATA(43) => X_Logic0_port, DATA(42) => X_Logic0_port, DATA(41) => 
               X_Logic0_port, DATA(40) => X_Logic0_port, 
         -- Connections to port 'DATA12'
         DATA(47) => X_Logic1_port, DATA(46) => X_Logic0_port, DATA(45) => 
               X_Logic0_port, DATA(44) => X_Logic0_port, 
         -- Connections to port 'DATA13'
         DATA(51) => X_Logic0_port, DATA(50) => X_Logic0_port, DATA(49) => 
               X_Logic0_port, DATA(48) => X_Logic0_port, 
         -- Connections to port 'DATA14'
         DATA(55) => X_Logic0_port, DATA(54) => X_Logic1_port, DATA(53) => 
               X_Logic1_port, DATA(52) => X_Logic1_port, 
         -- Connections to port 'DATA15'
         DATA(59) => X_Logic0_port, DATA(58) => X_Logic1_port, DATA(57) => 
               X_Logic1_port, DATA(56) => X_Logic1_port, 
         -- Connections to port 'DATA16'
         DATA(63) => X_Logic0_port, DATA(62) => X_Logic0_port, DATA(61) => 
               X_Logic0_port, DATA(60) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N48, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N49, 
         -- Connections to port 'CONTROL3'
         CONTROL(2) => N50, 
         -- Connections to port 'CONTROL4'
         CONTROL(3) => N51, 
         -- Connections to port 'CONTROL5'
         CONTROL(4) => N52, 
         -- Connections to port 'CONTROL6'
         CONTROL(5) => N53, 
         -- Connections to port 'CONTROL7'
         CONTROL(6) => N54, 
         -- Connections to port 'CONTROL8'
         CONTROL(7) => N55, 
         -- Connections to port 'CONTROL9'
         CONTROL(8) => N56, 
         -- Connections to port 'CONTROL10'
         CONTROL(9) => N57, 
         -- Connections to port 'CONTROL11'
         CONTROL(10) => N58, 
         -- Connections to port 'CONTROL12'
         CONTROL(11) => N59, 
         -- Connections to port 'CONTROL13'
         CONTROL(12) => N60, 
         -- Connections to port 'CONTROL14'
         CONTROL(13) => N61, 
         -- Connections to port 'CONTROL15'
         CONTROL(14) => N62, 
         -- Connections to port 'CONTROL16'
         CONTROL(15) => N63, 
         -- Connections to port 'Z'
         Z(3) => bdi_type_3_port, Z(2) => bdi_type_2_port, Z(1) => 
               bdi_type_1_port, Z(0) => bdi_type_0_port );
         X_Logic1_port <= '1';
         X_Logic0_port <= '0';
   B_64 : GTECH_BUF port map( A => N64, Z => last_flit_of_segment);
   C1063 : GTECH_OR2 port map( A => N97, B => N80, Z => N131);
   C1064 : GTECH_OR2 port map( A => N114, B => N131, Z => N132);
   C1065 : GTECH_OR2 port map( A => N130, B => N132, Z => N133);
   I_31 : GTECH_NOT port map( A => N133, Z => N134);
   C1071 : GTECH_OR2 port map( A => N166, B => N150, Z => N199);
   C1072 : GTECH_OR2 port map( A => N182, B => N199, Z => N200);
   C1073 : GTECH_OR2 port map( A => N198, B => N200, Z => N201);
   I_32 : GTECH_NOT port map( A => N201, Z => N202);
   I_33 : GTECH_NOT port map( A => sel_sdi_length, Z => N203);
   I_34 : GTECH_NOT port map( A => last_flit_of_segment, Z => N204);
   C1081 : GTECH_AND2 port map( A => eoi_flag, B => last_flit_of_segment, Z => 
                           bdi_eoi_internal);
   C1082 : GTECH_AND2 port map( A => eot_flag, B => last_flit_of_segment, Z => 
                           bdi_eot_internal);
   I_35 : GTECH_NOT port map( A => rst, Z => N205);
   I_36 : GTECH_NOT port map( A => pr_state_3_port, Z => N210);
   I_37 : GTECH_NOT port map( A => pr_state_2_port, Z => N211);
   I_38 : GTECH_NOT port map( A => pr_state_1_port, Z => N212);
   I_39 : GTECH_NOT port map( A => pr_state_0_port, Z => N213);
   I_40 : GTECH_NOT port map( A => N219, Z => N220);
   I_41 : GTECH_NOT port map( A => N223, Z => N224);
   I_42 : GTECH_NOT port map( A => N227, Z => N228);
   I_43 : GTECH_NOT port map( A => N231, Z => N232);
   I_44 : GTECH_NOT port map( A => N235, Z => N236);
   I_45 : GTECH_NOT port map( A => N239, Z => N240);
   I_46 : GTECH_NOT port map( A => N243, Z => N244);
   I_47 : GTECH_NOT port map( A => N247, Z => N248);
   I_48 : GTECH_NOT port map( A => N251, Z => N252);
   I_49 : GTECH_NOT port map( A => N255, Z => N256);
   I_50 : GTECH_NOT port map( A => N259, Z => N260);
   I_51 : GTECH_NOT port map( A => N263, Z => N264);
   I_52 : GTECH_NOT port map( A => N267, Z => N268);
   I_53 : GTECH_NOT port map( A => N271, Z => N272);
   C1150 : GTECH_AND2 port map( A => N527, B => cmd_ready_port, Z => N276);
   C1151 : GTECH_OR2 port map( A => N517, B => N521, Z => N527);
   I_54 : GTECH_NOT port map( A => N276, Z => N277);
   C1154 : GTECH_AND2 port map( A => N503, B => cmd_ready_port, Z => N278);
   I_55 : GTECH_NOT port map( A => sdi_valid_port, Z => N286);
   C1159 : GTECH_AND2 port map( A => N528, B => last_flit_of_segment, Z => N287
                           );
   C1160 : GTECH_AND2 port map( A => sdi_valid_port, B => key_ready_p, Z => 
                           N528);
   C1162 : GTECH_AND2 port map( A => N529, B => last_flit_of_segment, Z => N289
                           );
   C1163 : GTECH_AND2 port map( A => pdi_valid_port, B => bdi_ready_p, Z => 
                           N529);
   C1165 : GTECH_AND2 port map( A => N483, B => eot_flag, Z => N291);
   C1167 : GTECH_AND2 port map( A => N530, B => last_flit_of_segment, Z => N296
                           );
   C1168 : GTECH_AND2 port map( A => pdi_valid_port, B => bdi_ready_p, Z => 
                           N530);
   I_56 : GTECH_NOT port map( A => N296, Z => N297);
   I_57 : GTECH_NOT port map( A => eot_flag, Z => N298);
   C1174 : GTECH_AND2 port map( A => pdi_valid_port, B => cmd_ready_port, Z => 
                           N302);
   I_58 : GTECH_NOT port map( A => N302, Z => N303);
   C1177 : GTECH_AND2 port map( A => N499, B => eot_flag, Z => N304);
   I_59 : GTECH_NOT port map( A => N304, Z => N305);
   C1181 : GTECH_AND2 port map( A => N531, B => last_flit_of_segment, Z => N312
                           );
   C1182 : GTECH_AND2 port map( A => pdi_valid_port, B => bdi_ready_p, Z => 
                           N531);
   I_60 : GTECH_NOT port map( A => N312, Z => N313);
   C1189 : GTECH_AND2 port map( A => pdi_valid_port, B => last_flit_of_segment,
                           Z => N319);
   I_61 : GTECH_NOT port map( A => N319, Z => N320);
   C1193 : GTECH_AND2 port map( A => N532, B => last_flit_of_segment, Z => N324
                           );
   C1194 : GTECH_AND2 port map( A => pdi_valid_port, B => bdi_ready_p, Z => 
                           N532);
   I_62 : GTECH_NOT port map( A => N324, Z => N325);
   I_63 : GTECH_NOT port map( A => bdi_ready_p, Z => N328);
   I_64 : GTECH_NOT port map( A => N334, Z => N335);
   I_65 : GTECH_NOT port map( A => N338, Z => N339);
   I_66 : GTECH_NOT port map( A => N342, Z => N343);
   I_67 : GTECH_NOT port map( A => N346, Z => N347);
   I_68 : GTECH_NOT port map( A => N350, Z => N351);
   I_69 : GTECH_NOT port map( A => N354, Z => N355);
   I_70 : GTECH_NOT port map( A => N358, Z => N359);
   I_71 : GTECH_NOT port map( A => N362, Z => N363);
   I_72 : GTECH_NOT port map( A => N366, Z => N367);
   I_73 : GTECH_NOT port map( A => N370, Z => N371);
   I_74 : GTECH_NOT port map( A => N374, Z => N375);
   I_75 : GTECH_NOT port map( A => N378, Z => N379);
   I_76 : GTECH_NOT port map( A => N382, Z => N383);
   I_77 : GTECH_NOT port map( A => N386, Z => N387);
   C1263 : GTECH_OR2 port map( A => N508, B => N513, Z => N391);
   I_78 : GTECH_NOT port map( A => N391, Z => N392);
   I_79 : GTECH_NOT port map( A => pdi_valid_port, Z => N393);
   C1271 : GTECH_AND2 port map( A => sdi_valid_port, B => key_ready_p, Z => 
                           N402);
   C1272 : GTECH_AND2 port map( A => pdi_valid_port, B => bdi_ready_p, Z => 
                           N403);
   C1273 : GTECH_AND2 port map( A => pdi_valid_port, B => bdi_ready_p, Z => 
                           N404);
   C1275 : GTECH_AND2 port map( A => pdi_valid_port, B => bdi_ready_p, Z => 
                           N405);
   I_80 : GTECH_NOT port map( A => decrypt_port, Z => N406);
   C1279 : GTECH_AND2 port map( A => pdi_valid_port, B => bdi_ready_p, Z => 
                           N407);
   C1280 : GTECH_AND2 port map( A => pdi_valid_port, B => bdi_ready_p, Z => 
                           N411);
   C1281 : GTECH_OR2 port map( A => N335, B => N339, Z => N412);
   C1282 : GTECH_OR2 port map( A => N412, B => N343, Z => N413);
   C1283 : GTECH_OR2 port map( A => N413, B => N347, Z => N414);
   C1284 : GTECH_OR2 port map( A => N414, B => N351, Z => N415);
   C1285 : GTECH_OR2 port map( A => N415, B => N355, Z => N416);
   C1286 : GTECH_OR2 port map( A => N416, B => N359, Z => N417);
   C1287 : GTECH_OR2 port map( A => N417, B => N363, Z => N418);
   C1288 : GTECH_OR2 port map( A => N418, B => N367, Z => N419);
   C1289 : GTECH_OR2 port map( A => N419, B => N371, Z => N420);
   C1290 : GTECH_OR2 port map( A => N420, B => N375, Z => N421);
   C1291 : GTECH_OR2 port map( A => N421, B => N379, Z => N422);
   C1292 : GTECH_OR2 port map( A => N422, B => N383, Z => N423);
   C1293 : GTECH_OR2 port map( A => N423, B => N387, Z => N424);
   C1294 : GTECH_OR2 port map( A => N424, B => N390, Z => N425);
   I_81 : GTECH_NOT port map( A => N425, Z => N426);
   C1296 : GTECH_OR2 port map( A => N331, B => N335, Z => N427);
   C1297 : GTECH_OR2 port map( A => N427, B => N339, Z => N428);
   C1298 : GTECH_OR2 port map( A => N428, B => N343, Z => N429);
   C1299 : GTECH_AND2 port map( A => N393, B => N347, Z => N430);
   C1300 : GTECH_OR2 port map( A => N429, B => N430, Z => N431);
   C1301 : GTECH_OR2 port map( A => N431, B => N351, Z => N432);
   C1302 : GTECH_AND2 port map( A => N393, B => N355, Z => N433);
   C1303 : GTECH_OR2 port map( A => N432, B => N433, Z => N434);
   C1304 : GTECH_OR2 port map( A => N434, B => N359, Z => N435);
   C1305 : GTECH_AND2 port map( A => N303, B => N363, Z => N436);
   C1306 : GTECH_OR2 port map( A => N435, B => N436, Z => N437);
   C1307 : GTECH_OR2 port map( A => N437, B => N367, Z => N438);
   C1308 : GTECH_OR2 port map( A => N438, B => N371, Z => N439);
   C1309 : GTECH_OR2 port map( A => N439, B => N375, Z => N440);
   C1310 : GTECH_AND2 port map( A => N393, B => N379, Z => N441);
   C1311 : GTECH_OR2 port map( A => N440, B => N441, Z => N442);
   C1312 : GTECH_OR2 port map( A => N442, B => N383, Z => N443);
   C1313 : GTECH_OR2 port map( A => N443, B => N387, Z => N444);
   C1314 : GTECH_OR2 port map( A => N444, B => N390, Z => N445);
   I_82 : GTECH_NOT port map( A => N445, Z => N446);

end SYN_PreProcessor;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_LWC_1.all;

entity fwft_fifo_G_W32_G_LOG2DEPTH2 is

   port( clk, rst : in std_logic;  din : in std_logic_vector (31 downto 0);  
         din_valid : in std_logic;  din_ready : out std_logic;  dout : out 
         std_logic_vector (31 downto 0);  dout_valid : out std_logic;  
         dout_ready : in std_logic);

end fwft_fifo_G_W32_G_LOG2DEPTH2;

architecture SYN_structure of fwft_fifo_G_W32_G_LOG2DEPTH2 is

   component GTECH_AND2
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component GTECH_NOT
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component GTECH_OR2
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component GTECH_BUF
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX_OP
      generic( D0_width, D1_width, D2_width, D3_width, S0_width, S1_width, 
            Z_width : integer );
      port( D0 : in std_logic_vector(D0_width - 1 downto 0); D1 : in 
            std_logic_vector(D1_width - 1 downto 0); D2 : in 
            std_logic_vector(D2_width - 1 downto 0); D3 : in 
            std_logic_vector(D3_width - 1 downto 0); S0 : in 
            std_logic_vector(S0_width - 1 downto 0); S1 : in 
            std_logic_vector(S1_width - 1 downto 0); Z : out 
            std_logic_vector(Z_width - 1 downto 0) );
   end component;
   
   component SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
      generic ( ac_as_q, ac_as_qn, sc_ss_q : integer );
      port(
         clear, preset, enable, data_in, synch_clear, synch_preset, 
            synch_toggle, synch_enable, next_state, clocked_on : in std_logic;
         Q, QN : buffer std_logic
      );
   end component;
   
   signal N0, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, X_Logic1_port, 
      X_Logic0_port, clk_port, din_31_port, din_30_port, din_29_port, 
      din_28_port, din_27_port, din_26_port, din_25_port, din_24_port, 
      din_23_port, din_22_port, din_21_port, din_20_port, din_19_port, 
      din_18_port, din_17_port, din_16_port, din_15_port, din_14_port, 
      din_13_port, din_12_port, din_11_port, din_10_port, din_9_port, 
      din_8_port, din_7_port, din_6_port, din_5_port, din_4_port, din_3_port, 
      din_2_port, din_1_port, din_0_port, din_ready_port, dout_31_port, 
      dout_30_port, dout_29_port, dout_28_port, dout_27_port, dout_26_port, 
      dout_25_port, dout_24_port, dout_23_port, dout_22_port, dout_21_port, 
      dout_20_port, dout_19_port, dout_18_port, dout_17_port, dout_16_port, 
      dout_15_port, dout_14_port, dout_13_port, dout_12_port, dout_11_port, 
      dout_10_port, dout_9_port, dout_8_port, dout_7_port, dout_6_port, 
      dout_5_port, dout_4_port, dout_3_port, dout_2_port, dout_1_port, 
      dout_0_port, dout_valid_port, rd_ptr_s_1_port, rd_ptr_s_0_port, 
      mem_s_0_31_port, mem_s_0_30_port, mem_s_0_29_port, mem_s_0_28_port, 
      mem_s_0_27_port, mem_s_0_26_port, mem_s_0_25_port, mem_s_0_24_port, 
      mem_s_0_23_port, mem_s_0_22_port, mem_s_0_21_port, mem_s_0_20_port, 
      mem_s_0_19_port, mem_s_0_18_port, mem_s_0_17_port, mem_s_0_16_port, 
      mem_s_0_15_port, mem_s_0_14_port, mem_s_0_13_port, mem_s_0_12_port, 
      mem_s_0_11_port, mem_s_0_10_port, mem_s_0_9_port, mem_s_0_8_port, 
      mem_s_0_7_port, mem_s_0_6_port, mem_s_0_5_port, mem_s_0_4_port, 
      mem_s_0_3_port, mem_s_0_2_port, mem_s_0_1_port, mem_s_0_0_port, 
      mem_s_1_31_port, mem_s_1_30_port, mem_s_1_29_port, mem_s_1_28_port, 
      mem_s_1_27_port, mem_s_1_26_port, mem_s_1_25_port, mem_s_1_24_port, 
      mem_s_1_23_port, mem_s_1_22_port, mem_s_1_21_port, mem_s_1_20_port, 
      mem_s_1_19_port, mem_s_1_18_port, mem_s_1_17_port, mem_s_1_16_port, 
      mem_s_1_15_port, mem_s_1_14_port, mem_s_1_13_port, mem_s_1_12_port, 
      mem_s_1_11_port, mem_s_1_10_port, mem_s_1_9_port, mem_s_1_8_port, 
      mem_s_1_7_port, mem_s_1_6_port, mem_s_1_5_port, mem_s_1_4_port, 
      mem_s_1_3_port, mem_s_1_2_port, mem_s_1_1_port, mem_s_1_0_port, 
      mem_s_2_31_port, mem_s_2_30_port, mem_s_2_29_port, mem_s_2_28_port, 
      mem_s_2_27_port, mem_s_2_26_port, mem_s_2_25_port, mem_s_2_24_port, 
      mem_s_2_23_port, mem_s_2_22_port, mem_s_2_21_port, mem_s_2_20_port, 
      mem_s_2_19_port, mem_s_2_18_port, mem_s_2_17_port, mem_s_2_16_port, 
      mem_s_2_15_port, mem_s_2_14_port, mem_s_2_13_port, mem_s_2_12_port, 
      mem_s_2_11_port, mem_s_2_10_port, mem_s_2_9_port, mem_s_2_8_port, 
      mem_s_2_7_port, mem_s_2_6_port, mem_s_2_5_port, mem_s_2_4_port, 
      mem_s_2_3_port, mem_s_2_2_port, mem_s_2_1_port, mem_s_2_0_port, 
      mem_s_3_31_port, mem_s_3_30_port, mem_s_3_29_port, mem_s_3_28_port, 
      mem_s_3_27_port, mem_s_3_26_port, mem_s_3_25_port, mem_s_3_24_port, 
      mem_s_3_23_port, mem_s_3_22_port, mem_s_3_21_port, mem_s_3_20_port, 
      mem_s_3_19_port, mem_s_3_18_port, mem_s_3_17_port, mem_s_3_16_port, 
      mem_s_3_15_port, mem_s_3_14_port, mem_s_3_13_port, mem_s_3_12_port, 
      mem_s_3_11_port, mem_s_3_10_port, mem_s_3_9_port, mem_s_3_8_port, 
      mem_s_3_7_port, mem_s_3_6_port, mem_s_3_5_port, mem_s_3_4_port, 
      mem_s_3_3_port, mem_s_3_2_port, mem_s_3_1_port, mem_s_3_0_port, 
      entries_s_2_port, entries_s_1_port, entries_s_0_port, N12, full_s, N13, 
      empty_s, N14, wr_ptr_s_1_port, wr_ptr_s_0_port, N15, N16, N17, N18, N19, 
      N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34
      , N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, 
      N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63
      , N64, N65, N66, N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, n_1187
      , n_1188, n_1189, n_1190, n_1191, n_1192, n_1193, n_1194, n_1195, n_1196,
      n_1197, n_1198, n_1199, n_1200, n_1201, n_1202, n_1203, n_1204, n_1205, 
      n_1206, n_1207, n_1208, n_1209, n_1210, n_1211, n_1212, n_1213, n_1214, 
      n_1215, n_1216, n_1217, n_1218, n_1219, n_1220, n_1221, n_1222, n_1223, 
      n_1224, n_1225, n_1226, n_1227, n_1228, n_1229, n_1230, n_1231, n_1232, 
      n_1233, n_1234, n_1235, n_1236, n_1237, n_1238, n_1239, n_1240, n_1241, 
      n_1242, n_1243, n_1244, n_1245, n_1246, n_1247, n_1248, n_1249, n_1250, 
      n_1251, n_1252, n_1253, n_1254, n_1255, n_1256, n_1257, n_1258, n_1259, 
      n_1260, n_1261, n_1262, n_1263, n_1264, n_1265, n_1266, n_1267, n_1268, 
      n_1269, n_1270, n_1271, n_1272, n_1273, n_1274, n_1275, n_1276, n_1277, 
      n_1278, n_1279, n_1280, n_1281, n_1282, n_1283, n_1284, n_1285, n_1286, 
      n_1287, n_1288, n_1289, n_1290, n_1291, n_1292, n_1293, n_1294, n_1295, 
      n_1296, n_1297, n_1298, n_1299, n_1300, n_1301, n_1302, n_1303, n_1304, 
      n_1305, n_1306, n_1307, n_1308, n_1309, n_1310, n_1311, n_1312, n_1313, 
      n_1314, n_1315, n_1316, n_1317, n_1318, n_1319, n_1320, n_1321, n_1322, 
      n_1323, n_1324, n_1325 : std_logic;

begin
   clk_port <= clk;
   ( din_31_port, din_30_port, din_29_port, din_28_port, din_27_port, 
      din_26_port, din_25_port, din_24_port, din_23_port, din_22_port, 
      din_21_port, din_20_port, din_19_port, din_18_port, din_17_port, 
      din_16_port, din_15_port, din_14_port, din_13_port, din_12_port, 
      din_11_port, din_10_port, din_9_port, din_8_port, din_7_port, din_6_port,
      din_5_port, din_4_port, din_3_port, din_2_port, din_1_port, din_0_port ) 
      <= din;
   din_ready <= din_ready_port;
   dout <= ( dout_31_port, dout_30_port, dout_29_port, dout_28_port, 
      dout_27_port, dout_26_port, dout_25_port, dout_24_port, dout_23_port, 
      dout_22_port, dout_21_port, dout_20_port, dout_19_port, dout_18_port, 
      dout_17_port, dout_16_port, dout_15_port, dout_14_port, dout_13_port, 
      dout_12_port, dout_11_port, dout_10_port, dout_9_port, dout_8_port, 
      dout_7_port, dout_6_port, dout_5_port, dout_4_port, dout_3_port, 
      dout_2_port, dout_1_port, dout_0_port );
   dout_valid <= dout_valid_port;
   
   gte_77 : process ( X_Logic0_port, entries_s_2_port, entries_s_1_port, 
         entries_s_0_port, X_Logic1_port )
      variable A : SIGNED( 3 downto 0 );
      variable B : SIGNED( 3 downto 0 );
      variable Z : SIGNED( 0 downto 0 );
   begin
      A := ( X_Logic0_port, entries_s_2_port, entries_s_1_port, 
            entries_s_0_port );
      B := ( X_Logic0_port, X_Logic1_port, X_Logic0_port, X_Logic0_port );
      if ( A >= B ) then
         Z := ( others => '1' );
      else
         Z := ( others => '0' );
      end if;
      ( 0 => N12 ) <= Z;
   end process;
   
   lte_78 : process ( X_Logic0_port, entries_s_2_port, entries_s_1_port, 
         entries_s_0_port )
      variable A : SIGNED( 3 downto 0 );
      variable B : SIGNED( 0 downto 0 );
      variable Z : SIGNED( 0 downto 0 );
   begin
      A := ( X_Logic0_port, entries_s_2_port, entries_s_1_port, 
            entries_s_0_port );
      B := ( 0 => X_Logic0_port );
      if ( A <= B ) then
         Z := ( others => '1' );
      else
         Z := ( others => '0' );
      end if;
      ( 0 => N13 ) <= Z;
   end process;
   
   gte_107 : process ( X_Logic0_port, wr_ptr_s_1_port, wr_ptr_s_0_port, 
         X_Logic1_port )
      variable A : SIGNED( 2 downto 0 );
      variable B : SIGNED( 2 downto 0 );
      variable Z : SIGNED( 0 downto 0 );
   begin
      A := ( X_Logic0_port, wr_ptr_s_1_port, wr_ptr_s_0_port );
      B := ( X_Logic0_port, X_Logic1_port, X_Logic1_port );
      if ( A >= B ) then
         Z := ( others => '1' );
      else
         Z := ( others => '0' );
      end if;
      ( 0 => N37 ) <= Z;
   end process;
   
   gte_116 : process ( X_Logic0_port, rd_ptr_s_1_port, rd_ptr_s_0_port, 
         X_Logic1_port )
      variable A : SIGNED( 2 downto 0 );
      variable B : SIGNED( 2 downto 0 );
      variable Z : SIGNED( 0 downto 0 );
   begin
      A := ( X_Logic0_port, rd_ptr_s_1_port, rd_ptr_s_0_port );
      B := ( X_Logic0_port, X_Logic1_port, X_Logic1_port );
      if ( A >= B ) then
         Z := ( others => '1' );
      else
         Z := ( others => '0' );
      end if;
      ( 0 => N49 ) <= Z;
   end process;
   
   mem_s_reg_0_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N68, next_state => din_31_port, 
               clocked_on => clk_port, Q => mem_s_0_31_port, QN => n_1187);
   mem_s_reg_0_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N68, next_state => din_30_port, 
               clocked_on => clk_port, Q => mem_s_0_30_port, QN => n_1188);
   mem_s_reg_0_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N68, next_state => din_29_port, 
               clocked_on => clk_port, Q => mem_s_0_29_port, QN => n_1189);
   mem_s_reg_0_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N68, next_state => din_28_port, 
               clocked_on => clk_port, Q => mem_s_0_28_port, QN => n_1190);
   mem_s_reg_0_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N68, next_state => din_27_port, 
               clocked_on => clk_port, Q => mem_s_0_27_port, QN => n_1191);
   mem_s_reg_0_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N68, next_state => din_26_port, 
               clocked_on => clk_port, Q => mem_s_0_26_port, QN => n_1192);
   mem_s_reg_0_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N68, next_state => din_25_port, 
               clocked_on => clk_port, Q => mem_s_0_25_port, QN => n_1193);
   mem_s_reg_0_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N68, next_state => din_24_port, 
               clocked_on => clk_port, Q => mem_s_0_24_port, QN => n_1194);
   mem_s_reg_0_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N68, next_state => din_23_port, 
               clocked_on => clk_port, Q => mem_s_0_23_port, QN => n_1195);
   mem_s_reg_0_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N68, next_state => din_22_port, 
               clocked_on => clk_port, Q => mem_s_0_22_port, QN => n_1196);
   mem_s_reg_0_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N68, next_state => din_21_port, 
               clocked_on => clk_port, Q => mem_s_0_21_port, QN => n_1197);
   mem_s_reg_0_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N68, next_state => din_20_port, 
               clocked_on => clk_port, Q => mem_s_0_20_port, QN => n_1198);
   mem_s_reg_0_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N68, next_state => din_19_port, 
               clocked_on => clk_port, Q => mem_s_0_19_port, QN => n_1199);
   mem_s_reg_0_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N68, next_state => din_18_port, 
               clocked_on => clk_port, Q => mem_s_0_18_port, QN => n_1200);
   mem_s_reg_0_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N68, next_state => din_17_port, 
               clocked_on => clk_port, Q => mem_s_0_17_port, QN => n_1201);
   mem_s_reg_0_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N68, next_state => din_16_port, 
               clocked_on => clk_port, Q => mem_s_0_16_port, QN => n_1202);
   mem_s_reg_0_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N68, next_state => din_15_port, 
               clocked_on => clk_port, Q => mem_s_0_15_port, QN => n_1203);
   mem_s_reg_0_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N68, next_state => din_14_port, 
               clocked_on => clk_port, Q => mem_s_0_14_port, QN => n_1204);
   mem_s_reg_0_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N68, next_state => din_13_port, 
               clocked_on => clk_port, Q => mem_s_0_13_port, QN => n_1205);
   mem_s_reg_0_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N68, next_state => din_12_port, 
               clocked_on => clk_port, Q => mem_s_0_12_port, QN => n_1206);
   mem_s_reg_0_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N68, next_state => din_11_port, 
               clocked_on => clk_port, Q => mem_s_0_11_port, QN => n_1207);
   mem_s_reg_0_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N68, next_state => din_10_port, 
               clocked_on => clk_port, Q => mem_s_0_10_port, QN => n_1208);
   mem_s_reg_0_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N68, next_state => din_9_port, 
               clocked_on => clk_port, Q => mem_s_0_9_port, QN => n_1209);
   mem_s_reg_0_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N68, next_state => din_8_port, 
               clocked_on => clk_port, Q => mem_s_0_8_port, QN => n_1210);
   mem_s_reg_0_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N68, next_state => din_7_port, 
               clocked_on => clk_port, Q => mem_s_0_7_port, QN => n_1211);
   mem_s_reg_0_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N68, next_state => din_6_port, 
               clocked_on => clk_port, Q => mem_s_0_6_port, QN => n_1212);
   mem_s_reg_0_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N68, next_state => din_5_port, 
               clocked_on => clk_port, Q => mem_s_0_5_port, QN => n_1213);
   mem_s_reg_0_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N68, next_state => din_4_port, 
               clocked_on => clk_port, Q => mem_s_0_4_port, QN => n_1214);
   mem_s_reg_0_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N68, next_state => din_3_port, 
               clocked_on => clk_port, Q => mem_s_0_3_port, QN => n_1215);
   mem_s_reg_0_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N68, next_state => din_2_port, 
               clocked_on => clk_port, Q => mem_s_0_2_port, QN => n_1216);
   mem_s_reg_0_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N68, next_state => din_1_port, 
               clocked_on => clk_port, Q => mem_s_0_1_port, QN => n_1217);
   mem_s_reg_0_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N68, next_state => din_0_port, 
               clocked_on => clk_port, Q => mem_s_0_0_port, QN => n_1218);
   mem_s_reg_1_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N67, next_state => din_31_port, 
               clocked_on => clk_port, Q => mem_s_1_31_port, QN => n_1219);
   mem_s_reg_1_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N67, next_state => din_30_port, 
               clocked_on => clk_port, Q => mem_s_1_30_port, QN => n_1220);
   mem_s_reg_1_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N67, next_state => din_29_port, 
               clocked_on => clk_port, Q => mem_s_1_29_port, QN => n_1221);
   mem_s_reg_1_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N67, next_state => din_28_port, 
               clocked_on => clk_port, Q => mem_s_1_28_port, QN => n_1222);
   mem_s_reg_1_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N67, next_state => din_27_port, 
               clocked_on => clk_port, Q => mem_s_1_27_port, QN => n_1223);
   mem_s_reg_1_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N67, next_state => din_26_port, 
               clocked_on => clk_port, Q => mem_s_1_26_port, QN => n_1224);
   mem_s_reg_1_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N67, next_state => din_25_port, 
               clocked_on => clk_port, Q => mem_s_1_25_port, QN => n_1225);
   mem_s_reg_1_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N67, next_state => din_24_port, 
               clocked_on => clk_port, Q => mem_s_1_24_port, QN => n_1226);
   mem_s_reg_1_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N67, next_state => din_23_port, 
               clocked_on => clk_port, Q => mem_s_1_23_port, QN => n_1227);
   mem_s_reg_1_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N67, next_state => din_22_port, 
               clocked_on => clk_port, Q => mem_s_1_22_port, QN => n_1228);
   mem_s_reg_1_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N67, next_state => din_21_port, 
               clocked_on => clk_port, Q => mem_s_1_21_port, QN => n_1229);
   mem_s_reg_1_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N67, next_state => din_20_port, 
               clocked_on => clk_port, Q => mem_s_1_20_port, QN => n_1230);
   mem_s_reg_1_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N67, next_state => din_19_port, 
               clocked_on => clk_port, Q => mem_s_1_19_port, QN => n_1231);
   mem_s_reg_1_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N67, next_state => din_18_port, 
               clocked_on => clk_port, Q => mem_s_1_18_port, QN => n_1232);
   mem_s_reg_1_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N67, next_state => din_17_port, 
               clocked_on => clk_port, Q => mem_s_1_17_port, QN => n_1233);
   mem_s_reg_1_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N67, next_state => din_16_port, 
               clocked_on => clk_port, Q => mem_s_1_16_port, QN => n_1234);
   mem_s_reg_1_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N67, next_state => din_15_port, 
               clocked_on => clk_port, Q => mem_s_1_15_port, QN => n_1235);
   mem_s_reg_1_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N67, next_state => din_14_port, 
               clocked_on => clk_port, Q => mem_s_1_14_port, QN => n_1236);
   mem_s_reg_1_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N67, next_state => din_13_port, 
               clocked_on => clk_port, Q => mem_s_1_13_port, QN => n_1237);
   mem_s_reg_1_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N67, next_state => din_12_port, 
               clocked_on => clk_port, Q => mem_s_1_12_port, QN => n_1238);
   mem_s_reg_1_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N67, next_state => din_11_port, 
               clocked_on => clk_port, Q => mem_s_1_11_port, QN => n_1239);
   mem_s_reg_1_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N67, next_state => din_10_port, 
               clocked_on => clk_port, Q => mem_s_1_10_port, QN => n_1240);
   mem_s_reg_1_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N67, next_state => din_9_port, 
               clocked_on => clk_port, Q => mem_s_1_9_port, QN => n_1241);
   mem_s_reg_1_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N67, next_state => din_8_port, 
               clocked_on => clk_port, Q => mem_s_1_8_port, QN => n_1242);
   mem_s_reg_1_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N67, next_state => din_7_port, 
               clocked_on => clk_port, Q => mem_s_1_7_port, QN => n_1243);
   mem_s_reg_1_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N67, next_state => din_6_port, 
               clocked_on => clk_port, Q => mem_s_1_6_port, QN => n_1244);
   mem_s_reg_1_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N67, next_state => din_5_port, 
               clocked_on => clk_port, Q => mem_s_1_5_port, QN => n_1245);
   mem_s_reg_1_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N67, next_state => din_4_port, 
               clocked_on => clk_port, Q => mem_s_1_4_port, QN => n_1246);
   mem_s_reg_1_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N67, next_state => din_3_port, 
               clocked_on => clk_port, Q => mem_s_1_3_port, QN => n_1247);
   mem_s_reg_1_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N67, next_state => din_2_port, 
               clocked_on => clk_port, Q => mem_s_1_2_port, QN => n_1248);
   mem_s_reg_1_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N67, next_state => din_1_port, 
               clocked_on => clk_port, Q => mem_s_1_1_port, QN => n_1249);
   mem_s_reg_1_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N67, next_state => din_0_port, 
               clocked_on => clk_port, Q => mem_s_1_0_port, QN => n_1250);
   mem_s_reg_2_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N66, next_state => din_31_port, 
               clocked_on => clk_port, Q => mem_s_2_31_port, QN => n_1251);
   mem_s_reg_2_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N66, next_state => din_30_port, 
               clocked_on => clk_port, Q => mem_s_2_30_port, QN => n_1252);
   mem_s_reg_2_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N66, next_state => din_29_port, 
               clocked_on => clk_port, Q => mem_s_2_29_port, QN => n_1253);
   mem_s_reg_2_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N66, next_state => din_28_port, 
               clocked_on => clk_port, Q => mem_s_2_28_port, QN => n_1254);
   mem_s_reg_2_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N66, next_state => din_27_port, 
               clocked_on => clk_port, Q => mem_s_2_27_port, QN => n_1255);
   mem_s_reg_2_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N66, next_state => din_26_port, 
               clocked_on => clk_port, Q => mem_s_2_26_port, QN => n_1256);
   mem_s_reg_2_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N66, next_state => din_25_port, 
               clocked_on => clk_port, Q => mem_s_2_25_port, QN => n_1257);
   mem_s_reg_2_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N66, next_state => din_24_port, 
               clocked_on => clk_port, Q => mem_s_2_24_port, QN => n_1258);
   mem_s_reg_2_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N66, next_state => din_23_port, 
               clocked_on => clk_port, Q => mem_s_2_23_port, QN => n_1259);
   mem_s_reg_2_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N66, next_state => din_22_port, 
               clocked_on => clk_port, Q => mem_s_2_22_port, QN => n_1260);
   mem_s_reg_2_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N66, next_state => din_21_port, 
               clocked_on => clk_port, Q => mem_s_2_21_port, QN => n_1261);
   mem_s_reg_2_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N66, next_state => din_20_port, 
               clocked_on => clk_port, Q => mem_s_2_20_port, QN => n_1262);
   mem_s_reg_2_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N66, next_state => din_19_port, 
               clocked_on => clk_port, Q => mem_s_2_19_port, QN => n_1263);
   mem_s_reg_2_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N66, next_state => din_18_port, 
               clocked_on => clk_port, Q => mem_s_2_18_port, QN => n_1264);
   mem_s_reg_2_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N66, next_state => din_17_port, 
               clocked_on => clk_port, Q => mem_s_2_17_port, QN => n_1265);
   mem_s_reg_2_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N66, next_state => din_16_port, 
               clocked_on => clk_port, Q => mem_s_2_16_port, QN => n_1266);
   mem_s_reg_2_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N66, next_state => din_15_port, 
               clocked_on => clk_port, Q => mem_s_2_15_port, QN => n_1267);
   mem_s_reg_2_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N66, next_state => din_14_port, 
               clocked_on => clk_port, Q => mem_s_2_14_port, QN => n_1268);
   mem_s_reg_2_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N66, next_state => din_13_port, 
               clocked_on => clk_port, Q => mem_s_2_13_port, QN => n_1269);
   mem_s_reg_2_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N66, next_state => din_12_port, 
               clocked_on => clk_port, Q => mem_s_2_12_port, QN => n_1270);
   mem_s_reg_2_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N66, next_state => din_11_port, 
               clocked_on => clk_port, Q => mem_s_2_11_port, QN => n_1271);
   mem_s_reg_2_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N66, next_state => din_10_port, 
               clocked_on => clk_port, Q => mem_s_2_10_port, QN => n_1272);
   mem_s_reg_2_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N66, next_state => din_9_port, 
               clocked_on => clk_port, Q => mem_s_2_9_port, QN => n_1273);
   mem_s_reg_2_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N66, next_state => din_8_port, 
               clocked_on => clk_port, Q => mem_s_2_8_port, QN => n_1274);
   mem_s_reg_2_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N66, next_state => din_7_port, 
               clocked_on => clk_port, Q => mem_s_2_7_port, QN => n_1275);
   mem_s_reg_2_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N66, next_state => din_6_port, 
               clocked_on => clk_port, Q => mem_s_2_6_port, QN => n_1276);
   mem_s_reg_2_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N66, next_state => din_5_port, 
               clocked_on => clk_port, Q => mem_s_2_5_port, QN => n_1277);
   mem_s_reg_2_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N66, next_state => din_4_port, 
               clocked_on => clk_port, Q => mem_s_2_4_port, QN => n_1278);
   mem_s_reg_2_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N66, next_state => din_3_port, 
               clocked_on => clk_port, Q => mem_s_2_3_port, QN => n_1279);
   mem_s_reg_2_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N66, next_state => din_2_port, 
               clocked_on => clk_port, Q => mem_s_2_2_port, QN => n_1280);
   mem_s_reg_2_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N66, next_state => din_1_port, 
               clocked_on => clk_port, Q => mem_s_2_1_port, QN => n_1281);
   mem_s_reg_2_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N66, next_state => din_0_port, 
               clocked_on => clk_port, Q => mem_s_2_0_port, QN => n_1282);
   mem_s_reg_3_31_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N65, next_state => din_31_port, 
               clocked_on => clk_port, Q => mem_s_3_31_port, QN => n_1283);
   mem_s_reg_3_30_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N65, next_state => din_30_port, 
               clocked_on => clk_port, Q => mem_s_3_30_port, QN => n_1284);
   mem_s_reg_3_29_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N65, next_state => din_29_port, 
               clocked_on => clk_port, Q => mem_s_3_29_port, QN => n_1285);
   mem_s_reg_3_28_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N65, next_state => din_28_port, 
               clocked_on => clk_port, Q => mem_s_3_28_port, QN => n_1286);
   mem_s_reg_3_27_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N65, next_state => din_27_port, 
               clocked_on => clk_port, Q => mem_s_3_27_port, QN => n_1287);
   mem_s_reg_3_26_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N65, next_state => din_26_port, 
               clocked_on => clk_port, Q => mem_s_3_26_port, QN => n_1288);
   mem_s_reg_3_25_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N65, next_state => din_25_port, 
               clocked_on => clk_port, Q => mem_s_3_25_port, QN => n_1289);
   mem_s_reg_3_24_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N65, next_state => din_24_port, 
               clocked_on => clk_port, Q => mem_s_3_24_port, QN => n_1290);
   mem_s_reg_3_23_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N65, next_state => din_23_port, 
               clocked_on => clk_port, Q => mem_s_3_23_port, QN => n_1291);
   mem_s_reg_3_22_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N65, next_state => din_22_port, 
               clocked_on => clk_port, Q => mem_s_3_22_port, QN => n_1292);
   mem_s_reg_3_21_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N65, next_state => din_21_port, 
               clocked_on => clk_port, Q => mem_s_3_21_port, QN => n_1293);
   mem_s_reg_3_20_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N65, next_state => din_20_port, 
               clocked_on => clk_port, Q => mem_s_3_20_port, QN => n_1294);
   mem_s_reg_3_19_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N65, next_state => din_19_port, 
               clocked_on => clk_port, Q => mem_s_3_19_port, QN => n_1295);
   mem_s_reg_3_18_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N65, next_state => din_18_port, 
               clocked_on => clk_port, Q => mem_s_3_18_port, QN => n_1296);
   mem_s_reg_3_17_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N65, next_state => din_17_port, 
               clocked_on => clk_port, Q => mem_s_3_17_port, QN => n_1297);
   mem_s_reg_3_16_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N65, next_state => din_16_port, 
               clocked_on => clk_port, Q => mem_s_3_16_port, QN => n_1298);
   mem_s_reg_3_15_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N65, next_state => din_15_port, 
               clocked_on => clk_port, Q => mem_s_3_15_port, QN => n_1299);
   mem_s_reg_3_14_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N65, next_state => din_14_port, 
               clocked_on => clk_port, Q => mem_s_3_14_port, QN => n_1300);
   mem_s_reg_3_13_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N65, next_state => din_13_port, 
               clocked_on => clk_port, Q => mem_s_3_13_port, QN => n_1301);
   mem_s_reg_3_12_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N65, next_state => din_12_port, 
               clocked_on => clk_port, Q => mem_s_3_12_port, QN => n_1302);
   mem_s_reg_3_11_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N65, next_state => din_11_port, 
               clocked_on => clk_port, Q => mem_s_3_11_port, QN => n_1303);
   mem_s_reg_3_10_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N65, next_state => din_10_port, 
               clocked_on => clk_port, Q => mem_s_3_10_port, QN => n_1304);
   mem_s_reg_3_9_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N65, next_state => din_9_port, 
               clocked_on => clk_port, Q => mem_s_3_9_port, QN => n_1305);
   mem_s_reg_3_8_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N65, next_state => din_8_port, 
               clocked_on => clk_port, Q => mem_s_3_8_port, QN => n_1306);
   mem_s_reg_3_7_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N65, next_state => din_7_port, 
               clocked_on => clk_port, Q => mem_s_3_7_port, QN => n_1307);
   mem_s_reg_3_6_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N65, next_state => din_6_port, 
               clocked_on => clk_port, Q => mem_s_3_6_port, QN => n_1308);
   mem_s_reg_3_5_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N65, next_state => din_5_port, 
               clocked_on => clk_port, Q => mem_s_3_5_port, QN => n_1309);
   mem_s_reg_3_4_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N65, next_state => din_4_port, 
               clocked_on => clk_port, Q => mem_s_3_4_port, QN => n_1310);
   mem_s_reg_3_3_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N65, next_state => din_3_port, 
               clocked_on => clk_port, Q => mem_s_3_3_port, QN => n_1311);
   mem_s_reg_3_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N65, next_state => din_2_port, 
               clocked_on => clk_port, Q => mem_s_3_2_port, QN => n_1312);
   mem_s_reg_3_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N65, next_state => din_1_port, 
               clocked_on => clk_port, Q => mem_s_3_1_port, QN => n_1313);
   mem_s_reg_3_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N65, next_state => din_0_port, 
               clocked_on => clk_port, Q => mem_s_3_0_port, QN => n_1314);
   wr_ptr_s_reg_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N55, next_state => N57, 
               clocked_on => clk_port, Q => wr_ptr_s_1_port, QN => n_1315);
   wr_ptr_s_reg_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N55, next_state => N56, 
               clocked_on => clk_port, Q => wr_ptr_s_0_port, QN => n_1316);
   rd_ptr_s_reg_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N58, next_state => N60, 
               clocked_on => clk_port, Q => rd_ptr_s_1_port, QN => n_1317);
   rd_ptr_s_reg_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N58, next_state => N59, 
               clocked_on => clk_port, Q => rd_ptr_s_0_port, QN => n_1318);
   entries_s_reg_2_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N61, next_state => N64, 
               clocked_on => clk_port, Q => entries_s_2_port, QN => n_1319);
   entries_s_reg_1_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N61, next_state => N63, 
               clocked_on => clk_port, Q => entries_s_1_port, QN => n_1320);
   entries_s_reg_0_inst : SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT
         generic map ( ac_as_q => 5, ac_as_qn => 5, sc_ss_q => 5 )
         port map ( clear => X_Logic0_port, preset => X_Logic0_port, enable => 
               X_Logic0_port, data_in => X_Logic0_port, synch_clear => 
               X_Logic0_port, synch_preset => X_Logic0_port, synch_toggle => 
               X_Logic0_port, synch_enable => N61, next_state => N62, 
               clocked_on => clk_port, Q => entries_s_0_port, QN => n_1321);
   I_0 : GTECH_NOT port map( A => din_valid, Z => N69);
   I_1 : GTECH_NOT port map( A => din_ready_port, Z => N70);
   I_2 : GTECH_NOT port map( A => dout_valid_port, Z => N71);
   I_3 : GTECH_NOT port map( A => dout_ready, Z => N72);
   add_98 : process ( entries_s_2_port, entries_s_1_port, entries_s_0_port, 
         X_Logic0_port, X_Logic1_port )
      variable A : SIGNED( 2 downto 0 );
      variable B : SIGNED( 2 downto 0 );
      variable Z : SIGNED( 2 downto 0 );
   begin
      A := ( entries_s_2_port, entries_s_1_port, entries_s_0_port );
      B := ( X_Logic0_port, X_Logic0_port, X_Logic1_port );
      Z := A + B;
      ( N20, N19, N18 ) <= Z;
   end process;
   
   sub_101 : process ( entries_s_2_port, entries_s_1_port, entries_s_0_port, 
         X_Logic0_port, X_Logic1_port )
      variable A : SIGNED( 2 downto 0 );
      variable B : SIGNED( 2 downto 0 );
      variable Z : SIGNED( 2 downto 0 );
   begin
      A := ( entries_s_2_port, entries_s_1_port, entries_s_0_port );
      B := ( X_Logic0_port, X_Logic0_port, X_Logic1_port );
      Z := A - B;
      ( N25, N24, N23 ) <= Z;
   end process;
   
   add_110 : process ( wr_ptr_s_1_port, wr_ptr_s_0_port, X_Logic0_port, 
         X_Logic1_port )
      variable A : SIGNED( 1 downto 0 );
      variable B : SIGNED( 1 downto 0 );
      variable Z : SIGNED( 1 downto 0 );
   begin
      A := ( wr_ptr_s_1_port, wr_ptr_s_0_port );
      B := ( X_Logic0_port, X_Logic1_port );
      Z := A + B;
      ( N40, N39 ) <= Z;
   end process;
   
   add_119 : process ( rd_ptr_s_1_port, rd_ptr_s_0_port, X_Logic0_port, 
         X_Logic1_port )
      variable A : SIGNED( 1 downto 0 );
      variable B : SIGNED( 1 downto 0 );
      variable Z : SIGNED( 1 downto 0 );
   begin
      A := ( rd_ptr_s_1_port, rd_ptr_s_0_port );
      B := ( X_Logic0_port, X_Logic1_port );
      Z := A + B;
      ( N52, N51 ) <= Z;
   end process;
   
   C635 : GTECH_AND2 port map( A => wr_ptr_s_0_port, B => wr_ptr_s_1_port, Z =>
                           N36);
   C636 : GTECH_AND2 port map( A => N0, B => wr_ptr_s_1_port, Z => N35);
   I_4 : GTECH_NOT port map( A => wr_ptr_s_0_port, Z => N0);
   C637 : GTECH_AND2 port map( A => wr_ptr_s_0_port, B => N1, Z => N34);
   I_5 : GTECH_NOT port map( A => wr_ptr_s_1_port, Z => N1);
   C638 : GTECH_AND2 port map( A => N2, B => N3, Z => N33);
   I_6 : GTECH_NOT port map( A => wr_ptr_s_0_port, Z => N2);
   I_7 : GTECH_NOT port map( A => wr_ptr_s_1_port, Z => N3);
   C639_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic1_port, 
         -- Connections to port 'DATA2'
         DATA(1) => N22, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N4, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N17, 
         -- Connections to port 'Z'
         Z(0) => N26 );
   B_0 : GTECH_BUF port map( A => N16, Z => N4);
   C640_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 3 )
      port map(
         -- Connections to port 'DATA1'
         DATA(2) => N20, DATA(1) => N19, DATA(0) => N18, 
         -- Connections to port 'DATA2'
         DATA(5) => N25, DATA(4) => N24, DATA(3) => N23, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N4, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N17, 
         -- Connections to port 'Z'
         Z(2) => N29, Z(1) => N28, Z(0) => N27 );
   C641_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 2 )
      port map(
         -- Connections to port 'DATA1'
         DATA(1) => X_Logic0_port, DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(3) => N40, DATA(2) => N39, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N5, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N38, 
         -- Connections to port 'Z'
         Z(1) => N42, Z(0) => N41 );
   B_1 : GTECH_BUF port map( A => N37, Z => N5);
   C642_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 4 )
      port map(
         -- Connections to port 'DATA1'
         DATA(3) => N33, DATA(2) => N34, DATA(1) => N35, DATA(0) => N36, 
         -- Connections to port 'DATA2'
         DATA(7) => X_Logic0_port, DATA(6) => X_Logic0_port, DATA(5) => 
               X_Logic0_port, DATA(4) => X_Logic0_port, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N6, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N31, 
         -- Connections to port 'Z'
         Z(3) => N46, Z(2) => N45, Z(1) => N44, Z(0) => N43 );
   B_2 : GTECH_BUF port map( A => N30, Z => N6);
   C643_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 2 )
      port map(
         -- Connections to port 'DATA1'
         DATA(1) => X_Logic0_port, DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(3) => N52, DATA(2) => N51, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N7, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N50, 
         -- Connections to port 'Z'
         Z(1) => N54, Z(0) => N53 );
   B_3 : GTECH_BUF port map( A => N49, Z => N7);
   C644_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic1_port, 
         -- Connections to port 'DATA2'
         DATA(1) => N30, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N8, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N9, 
         -- Connections to port 'Z'
         Z(0) => N55 );
   B_4 : GTECH_BUF port map( A => rst, Z => N8);
   B_5 : GTECH_BUF port map( A => N14, Z => N9);
   C645_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 2 )
      port map(
         -- Connections to port 'DATA1'
         DATA(1) => X_Logic0_port, DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(3) => N42, DATA(2) => N41, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N8, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N9, 
         -- Connections to port 'Z'
         Z(1) => N57, Z(0) => N56 );
   C646_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic1_port, 
         -- Connections to port 'DATA2'
         DATA(1) => N47, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N8, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N9, 
         -- Connections to port 'Z'
         Z(0) => N58 );
   C647_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 2 )
      port map(
         -- Connections to port 'DATA1'
         DATA(1) => X_Logic0_port, DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(3) => N54, DATA(2) => N53, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N8, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N9, 
         -- Connections to port 'Z'
         Z(1) => N60, Z(0) => N59 );
   C648_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 1 )
      port map(
         -- Connections to port 'DATA1'
         DATA(0) => X_Logic1_port, 
         -- Connections to port 'DATA2'
         DATA(1) => N26, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N8, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N9, 
         -- Connections to port 'Z'
         Z(0) => N61 );
   C649_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 3 )
      port map(
         -- Connections to port 'DATA1'
         DATA(2) => X_Logic0_port, DATA(1) => X_Logic0_port, DATA(0) => 
               X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(5) => N29, DATA(4) => N28, DATA(3) => N27, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N8, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N9, 
         -- Connections to port 'Z'
         Z(2) => N64, Z(1) => N63, Z(0) => N62 );
   C650_cell : SELECT_OP
      generic map ( num_inputs => 2, input_width => 4 )
      port map(
         -- Connections to port 'DATA1'
         DATA(3) => X_Logic0_port, DATA(2) => X_Logic0_port, DATA(1) => 
               X_Logic0_port, DATA(0) => X_Logic0_port, 
         -- Connections to port 'DATA2'
         DATA(7) => N46, DATA(6) => N45, DATA(5) => N44, DATA(4) => N43, 
         -- Connections to port 'CONTROL1'
         CONTROL(0) => N8, 
         -- Connections to port 'CONTROL2'
         CONTROL(1) => N9, 
         -- Connections to port 'Z'
         Z(3) => N68, Z(2) => N67, Z(1) => N66, Z(0) => N65 );
   C651 : MUX_OP
      generic map ( D0_width => 32, D1_width => 32, D2_width => 32, D3_width =>
            32, S0_width => 1, S1_width => 1, Z_width => 32 )
      port map(
         -- Connections to port 'D0'
         D0(31) => mem_s_0_0_port, D0(30) => mem_s_0_1_port, D0(29) => 
               mem_s_0_2_port, D0(28) => mem_s_0_3_port, D0(27) => 
               mem_s_0_4_port, D0(26) => mem_s_0_5_port, D0(25) => 
               mem_s_0_6_port, D0(24) => mem_s_0_7_port, D0(23) => 
               mem_s_0_8_port, D0(22) => mem_s_0_9_port, D0(21) => 
               mem_s_0_10_port, D0(20) => mem_s_0_11_port, D0(19) => 
               mem_s_0_12_port, D0(18) => mem_s_0_13_port, D0(17) => 
               mem_s_0_14_port, D0(16) => mem_s_0_15_port, D0(15) => 
               mem_s_0_16_port, D0(14) => mem_s_0_17_port, D0(13) => 
               mem_s_0_18_port, D0(12) => mem_s_0_19_port, D0(11) => 
               mem_s_0_20_port, D0(10) => mem_s_0_21_port, D0(9) => 
               mem_s_0_22_port, D0(8) => mem_s_0_23_port, D0(7) => 
               mem_s_0_24_port, D0(6) => mem_s_0_25_port, D0(5) => 
               mem_s_0_26_port, D0(4) => mem_s_0_27_port, D0(3) => 
               mem_s_0_28_port, D0(2) => mem_s_0_29_port, D0(1) => 
               mem_s_0_30_port, D0(0) => mem_s_0_31_port, 
         -- Connections to port 'D1'
         D1(31) => mem_s_1_0_port, D1(30) => mem_s_1_1_port, D1(29) => 
               mem_s_1_2_port, D1(28) => mem_s_1_3_port, D1(27) => 
               mem_s_1_4_port, D1(26) => mem_s_1_5_port, D1(25) => 
               mem_s_1_6_port, D1(24) => mem_s_1_7_port, D1(23) => 
               mem_s_1_8_port, D1(22) => mem_s_1_9_port, D1(21) => 
               mem_s_1_10_port, D1(20) => mem_s_1_11_port, D1(19) => 
               mem_s_1_12_port, D1(18) => mem_s_1_13_port, D1(17) => 
               mem_s_1_14_port, D1(16) => mem_s_1_15_port, D1(15) => 
               mem_s_1_16_port, D1(14) => mem_s_1_17_port, D1(13) => 
               mem_s_1_18_port, D1(12) => mem_s_1_19_port, D1(11) => 
               mem_s_1_20_port, D1(10) => mem_s_1_21_port, D1(9) => 
               mem_s_1_22_port, D1(8) => mem_s_1_23_port, D1(7) => 
               mem_s_1_24_port, D1(6) => mem_s_1_25_port, D1(5) => 
               mem_s_1_26_port, D1(4) => mem_s_1_27_port, D1(3) => 
               mem_s_1_28_port, D1(2) => mem_s_1_29_port, D1(1) => 
               mem_s_1_30_port, D1(0) => mem_s_1_31_port, 
         -- Connections to port 'D2'
         D2(31) => mem_s_2_0_port, D2(30) => mem_s_2_1_port, D2(29) => 
               mem_s_2_2_port, D2(28) => mem_s_2_3_port, D2(27) => 
               mem_s_2_4_port, D2(26) => mem_s_2_5_port, D2(25) => 
               mem_s_2_6_port, D2(24) => mem_s_2_7_port, D2(23) => 
               mem_s_2_8_port, D2(22) => mem_s_2_9_port, D2(21) => 
               mem_s_2_10_port, D2(20) => mem_s_2_11_port, D2(19) => 
               mem_s_2_12_port, D2(18) => mem_s_2_13_port, D2(17) => 
               mem_s_2_14_port, D2(16) => mem_s_2_15_port, D2(15) => 
               mem_s_2_16_port, D2(14) => mem_s_2_17_port, D2(13) => 
               mem_s_2_18_port, D2(12) => mem_s_2_19_port, D2(11) => 
               mem_s_2_20_port, D2(10) => mem_s_2_21_port, D2(9) => 
               mem_s_2_22_port, D2(8) => mem_s_2_23_port, D2(7) => 
               mem_s_2_24_port, D2(6) => mem_s_2_25_port, D2(5) => 
               mem_s_2_26_port, D2(4) => mem_s_2_27_port, D2(3) => 
               mem_s_2_28_port, D2(2) => mem_s_2_29_port, D2(1) => 
               mem_s_2_30_port, D2(0) => mem_s_2_31_port, 
         -- Connections to port 'D3'
         D3(31) => mem_s_3_0_port, D3(30) => mem_s_3_1_port, D3(29) => 
               mem_s_3_2_port, D3(28) => mem_s_3_3_port, D3(27) => 
               mem_s_3_4_port, D3(26) => mem_s_3_5_port, D3(25) => 
               mem_s_3_6_port, D3(24) => mem_s_3_7_port, D3(23) => 
               mem_s_3_8_port, D3(22) => mem_s_3_9_port, D3(21) => 
               mem_s_3_10_port, D3(20) => mem_s_3_11_port, D3(19) => 
               mem_s_3_12_port, D3(18) => mem_s_3_13_port, D3(17) => 
               mem_s_3_14_port, D3(16) => mem_s_3_15_port, D3(15) => 
               mem_s_3_16_port, D3(14) => mem_s_3_17_port, D3(13) => 
               mem_s_3_18_port, D3(12) => mem_s_3_19_port, D3(11) => 
               mem_s_3_20_port, D3(10) => mem_s_3_21_port, D3(9) => 
               mem_s_3_22_port, D3(8) => mem_s_3_23_port, D3(7) => 
               mem_s_3_24_port, D3(6) => mem_s_3_25_port, D3(5) => 
               mem_s_3_26_port, D3(4) => mem_s_3_27_port, D3(3) => 
               mem_s_3_28_port, D3(2) => mem_s_3_29_port, D3(1) => 
               mem_s_3_30_port, D3(0) => mem_s_3_31_port, 
         -- Connections to port 'S0'
         S0(0) => N10, 
         -- Connections to port 'S1'
         S1(0) => N11, 
         -- Connections to port 'Z'
         Z(31) => dout_0_port, Z(30) => dout_1_port, Z(29) => dout_2_port, 
               Z(28) => dout_3_port, Z(27) => dout_4_port, Z(26) => dout_5_port
               , Z(25) => dout_6_port, Z(24) => dout_7_port, Z(23) => 
               dout_8_port, Z(22) => dout_9_port, Z(21) => dout_10_port, Z(20) 
               => dout_11_port, Z(19) => dout_12_port, Z(18) => dout_13_port, 
               Z(17) => dout_14_port, Z(16) => dout_15_port, Z(15) => 
               dout_16_port, Z(14) => dout_17_port, Z(13) => dout_18_port, 
               Z(12) => dout_19_port, Z(11) => dout_20_port, Z(10) => 
               dout_21_port, Z(9) => dout_22_port, Z(8) => dout_23_port, Z(7) 
               => dout_24_port, Z(6) => dout_25_port, Z(5) => dout_26_port, 
               Z(4) => dout_27_port, Z(3) => dout_28_port, Z(2) => dout_29_port
               , Z(1) => dout_30_port, Z(0) => dout_31_port
      );
   B_6 : GTECH_BUF port map( A => rd_ptr_s_0_port, Z => N10);
   B_7 : GTECH_BUF port map( A => rd_ptr_s_1_port, Z => N11);
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   B_8 : GTECH_BUF port map( A => N12, Z => full_s);
   B_9 : GTECH_BUF port map( A => N13, Z => empty_s);
   I_8 : GTECH_NOT port map( A => full_s, Z => din_ready_port);
   I_9 : GTECH_NOT port map( A => empty_s, Z => dout_valid_port);
   I_10 : GTECH_NOT port map( A => rst, Z => N14);
   B_10 : GTECH_BUF port map( A => N14, Z => N15);
   C662 : GTECH_AND2 port map( A => N73, B => N74, Z => N16);
   C663 : GTECH_AND2 port map( A => din_valid, B => din_ready_port, Z => N73);
   C664 : GTECH_OR2 port map( A => N71, B => N72, Z => N74);
   I_11 : GTECH_NOT port map( A => N16, Z => N17);
   C667 : GTECH_AND2 port map( A => N15, B => N16, Z => n_1322);
   C668 : GTECH_AND2 port map( A => N15, B => N17, Z => N21);
   C669 : GTECH_AND2 port map( A => N76, B => dout_ready, Z => N22);
   C670 : GTECH_AND2 port map( A => N75, B => dout_valid_port, Z => N76);
   C671 : GTECH_OR2 port map( A => N69, B => N70, Z => N75);
   C673 : GTECH_AND2 port map( A => N21, B => N22, Z => n_1323);
   C674 : GTECH_AND2 port map( A => din_valid, B => din_ready_port, Z => N30);
   I_12 : GTECH_NOT port map( A => N30, Z => N31);
   C677 : GTECH_AND2 port map( A => N15, B => N30, Z => N32);
   I_13 : GTECH_NOT port map( A => N37, Z => N38);
   C680 : GTECH_AND2 port map( A => N32, B => N38, Z => n_1324);
   C681 : GTECH_AND2 port map( A => dout_valid_port, B => dout_ready, Z => N47)
                           ;
   C683 : GTECH_AND2 port map( A => N15, B => N47, Z => N48);
   I_14 : GTECH_NOT port map( A => N49, Z => N50);
   C686 : GTECH_AND2 port map( A => N48, B => N50, Z => n_1325);

end SYN_structure;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_LWC_1.all;

entity LWC_1 is

   port( clk, rst : in std_logic;  pdi_data : in std_logic_vector (31 downto 0)
         ;  pdi_valid : in std_logic;  pdi_ready : out std_logic;  sdi_data : 
         in std_logic_vector (31 downto 0);  sdi_valid : in std_logic;  
         sdi_ready : out std_logic;  do_data : out std_logic_vector (31 downto 
         0);  do_ready : in std_logic;  do_valid, do_last : out std_logic);

end LWC_1;

architecture SYN_structure of LWC_1 is

   component fwft_fifo_G_W32_G_LOG2DEPTH2
      port( clk, rst : in std_logic;  din : in std_logic_vector (31 downto 0); 
            din_valid : in std_logic;  din_ready : out std_logic;  dout : out 
            std_logic_vector (31 downto 0);  dout_valid : out std_logic;  
            dout_ready : in std_logic);
   end component;
   
   component PostProcessor_2
      port( clk, rst : in std_logic;  bdo : in std_logic_vector (31 downto 0); 
            bdo_valid : in std_logic;  bdo_ready : out std_logic;  end_of_block
            : in std_logic;  bdo_type, bdo_valid_bytes : in std_logic_vector (3
            downto 0);  msg_auth : in std_logic;  msg_auth_ready : out 
            std_logic;  msg_auth_valid : in std_logic;  cmd : in 
            std_logic_vector (31 downto 0);  cmd_valid : in std_logic;  
            cmd_ready : out std_logic;  do_data : out std_logic_vector (31 
            downto 0);  do_valid, do_last : out std_logic;  do_ready : in 
            std_logic);
   end component;
   
   component CryptoCore_2
      port( clk, rst : in std_logic;  key : in std_logic_vector (31 downto 0); 
            key_valid : in std_logic;  key_ready : out std_logic;  bdi : in 
            std_logic_vector (31 downto 0);  bdi_valid : in std_logic;  
            bdi_ready : out std_logic;  bdi_pad_loc, bdi_valid_bytes : in 
            std_logic_vector (3 downto 0);  bdi_size : in std_logic_vector (2 
            downto 0);  bdi_eot, bdi_eoi : in std_logic;  bdi_type : in 
            std_logic_vector (3 downto 0);  decrypt_in, key_update, hash_in : 
            in std_logic;  bdo : out std_logic_vector (31 downto 0);  bdo_valid
            : out std_logic;  bdo_ready : in std_logic;  bdo_type, 
            bdo_valid_bytes : out std_logic_vector (3 downto 0);  end_of_block,
            msg_auth_valid : out std_logic;  msg_auth_ready : in std_logic;  
            msg_auth : out std_logic);
   end component;
   
   component PreProcessor_2
      port( clk, rst : in std_logic;  pdi_data : in std_logic_vector (31 downto
            0);  pdi_valid : in std_logic;  pdi_ready : out std_logic;  
            sdi_data : in std_logic_vector (31 downto 0);  sdi_valid : in 
            std_logic;  sdi_ready : out std_logic;  key : out std_logic_vector 
            (31 downto 0);  key_valid : out std_logic;  key_ready : in 
            std_logic;  bdi : out std_logic_vector (31 downto 0);  bdi_valid : 
            out std_logic;  bdi_ready : in std_logic;  bdi_pad_loc, 
            bdi_valid_bytes : out std_logic_vector (3 downto 0);  bdi_size : 
            out std_logic_vector (2 downto 0);  bdi_eot, bdi_eoi : out 
            std_logic;  bdi_type : out std_logic_vector (3 downto 0);  decrypt,
            hash, key_update : out std_logic;  cmd : out std_logic_vector (31 
            downto 0);  cmd_valid : out std_logic;  cmd_ready : in std_logic);
   end component;
   
   signal key_cipher_in_31_port, key_cipher_in_30_port, key_cipher_in_29_port, 
      key_cipher_in_28_port, key_cipher_in_27_port, key_cipher_in_26_port, 
      key_cipher_in_25_port, key_cipher_in_24_port, key_cipher_in_23_port, 
      key_cipher_in_22_port, key_cipher_in_21_port, key_cipher_in_20_port, 
      key_cipher_in_19_port, key_cipher_in_18_port, key_cipher_in_17_port, 
      key_cipher_in_16_port, key_cipher_in_15_port, key_cipher_in_14_port, 
      key_cipher_in_13_port, key_cipher_in_12_port, key_cipher_in_11_port, 
      key_cipher_in_10_port, key_cipher_in_9_port, key_cipher_in_8_port, 
      key_cipher_in_7_port, key_cipher_in_6_port, key_cipher_in_5_port, 
      key_cipher_in_4_port, key_cipher_in_3_port, key_cipher_in_2_port, 
      key_cipher_in_1_port, key_cipher_in_0_port, key_valid_cipher_in, 
      key_ready_cipher_in, bdi_cipher_in_31_port, bdi_cipher_in_30_port, 
      bdi_cipher_in_29_port, bdi_cipher_in_28_port, bdi_cipher_in_27_port, 
      bdi_cipher_in_26_port, bdi_cipher_in_25_port, bdi_cipher_in_24_port, 
      bdi_cipher_in_23_port, bdi_cipher_in_22_port, bdi_cipher_in_21_port, 
      bdi_cipher_in_20_port, bdi_cipher_in_19_port, bdi_cipher_in_18_port, 
      bdi_cipher_in_17_port, bdi_cipher_in_16_port, bdi_cipher_in_15_port, 
      bdi_cipher_in_14_port, bdi_cipher_in_13_port, bdi_cipher_in_12_port, 
      bdi_cipher_in_11_port, bdi_cipher_in_10_port, bdi_cipher_in_9_port, 
      bdi_cipher_in_8_port, bdi_cipher_in_7_port, bdi_cipher_in_6_port, 
      bdi_cipher_in_5_port, bdi_cipher_in_4_port, bdi_cipher_in_3_port, 
      bdi_cipher_in_2_port, bdi_cipher_in_1_port, bdi_cipher_in_0_port, 
      bdi_valid_cipher_in, bdi_ready_cipher_in, bdi_pad_loc_cipher_in_3_port, 
      bdi_pad_loc_cipher_in_2_port, bdi_pad_loc_cipher_in_1_port, 
      bdi_pad_loc_cipher_in_0_port, bdi_valid_bytes_cipher_in_3_port, 
      bdi_valid_bytes_cipher_in_2_port, bdi_valid_bytes_cipher_in_1_port, 
      bdi_valid_bytes_cipher_in_0_port, bdi_size_cipher_in_2_port, 
      bdi_size_cipher_in_1_port, bdi_size_cipher_in_0_port, bdi_eot_cipher_in, 
      bdi_eoi_cipher_in, bdi_type_cipher_in_3_port, bdi_type_cipher_in_2_port, 
      bdi_type_cipher_in_1_port, bdi_type_cipher_in_0_port, decrypt_cipher_in, 
      hash_cipher_in, key_update_cipher_in, cmd_FIFO_in_31_port, 
      cmd_FIFO_in_30_port, cmd_FIFO_in_29_port, cmd_FIFO_in_28_port, 
      cmd_FIFO_in_27_port, cmd_FIFO_in_26_port, cmd_FIFO_in_25_port, 
      cmd_FIFO_in_24_port, cmd_FIFO_in_23_port, cmd_FIFO_in_22_port, 
      cmd_FIFO_in_21_port, cmd_FIFO_in_20_port, cmd_FIFO_in_19_port, 
      cmd_FIFO_in_18_port, cmd_FIFO_in_17_port, cmd_FIFO_in_16_port, 
      cmd_FIFO_in_15_port, cmd_FIFO_in_14_port, cmd_FIFO_in_13_port, 
      cmd_FIFO_in_12_port, cmd_FIFO_in_11_port, cmd_FIFO_in_10_port, 
      cmd_FIFO_in_9_port, cmd_FIFO_in_8_port, cmd_FIFO_in_7_port, 
      cmd_FIFO_in_6_port, cmd_FIFO_in_5_port, cmd_FIFO_in_4_port, 
      cmd_FIFO_in_3_port, cmd_FIFO_in_2_port, cmd_FIFO_in_1_port, 
      cmd_FIFO_in_0_port, cmd_valid_FIFO_in, cmd_ready_FIFO_in, 
      bdo_cipher_out_31_port, bdo_cipher_out_30_port, bdo_cipher_out_29_port, 
      bdo_cipher_out_28_port, bdo_cipher_out_27_port, bdo_cipher_out_26_port, 
      bdo_cipher_out_25_port, bdo_cipher_out_24_port, bdo_cipher_out_23_port, 
      bdo_cipher_out_22_port, bdo_cipher_out_21_port, bdo_cipher_out_20_port, 
      bdo_cipher_out_19_port, bdo_cipher_out_18_port, bdo_cipher_out_17_port, 
      bdo_cipher_out_16_port, bdo_cipher_out_15_port, bdo_cipher_out_14_port, 
      bdo_cipher_out_13_port, bdo_cipher_out_12_port, bdo_cipher_out_11_port, 
      bdo_cipher_out_10_port, bdo_cipher_out_9_port, bdo_cipher_out_8_port, 
      bdo_cipher_out_7_port, bdo_cipher_out_6_port, bdo_cipher_out_5_port, 
      bdo_cipher_out_4_port, bdo_cipher_out_3_port, bdo_cipher_out_2_port, 
      bdo_cipher_out_1_port, bdo_cipher_out_0_port, bdo_valid_cipher_out, 
      bdo_ready_cipher_out, bdo_type_cipher_out_3_port, 
      bdo_type_cipher_out_2_port, bdo_type_cipher_out_1_port, 
      bdo_type_cipher_out_0_port, bdo_valid_bytes_cipher_out_3_port, 
      bdo_valid_bytes_cipher_out_2_port, bdo_valid_bytes_cipher_out_1_port, 
      bdo_valid_bytes_cipher_out_0_port, end_of_block_cipher_out, 
      msg_auth_valid, msg_auth_ready, msg_auth, cmd_FIFO_out_31_port, 
      cmd_FIFO_out_30_port, cmd_FIFO_out_29_port, cmd_FIFO_out_28_port, 
      cmd_FIFO_out_27_port, cmd_FIFO_out_26_port, cmd_FIFO_out_25_port, 
      cmd_FIFO_out_24_port, cmd_FIFO_out_23_port, cmd_FIFO_out_22_port, 
      cmd_FIFO_out_21_port, cmd_FIFO_out_20_port, cmd_FIFO_out_19_port, 
      cmd_FIFO_out_18_port, cmd_FIFO_out_17_port, cmd_FIFO_out_16_port, 
      cmd_FIFO_out_15_port, cmd_FIFO_out_14_port, cmd_FIFO_out_13_port, 
      cmd_FIFO_out_12_port, cmd_FIFO_out_11_port, cmd_FIFO_out_10_port, 
      cmd_FIFO_out_9_port, cmd_FIFO_out_8_port, cmd_FIFO_out_7_port, 
      cmd_FIFO_out_6_port, cmd_FIFO_out_5_port, cmd_FIFO_out_4_port, 
      cmd_FIFO_out_3_port, cmd_FIFO_out_2_port, cmd_FIFO_out_1_port, 
      cmd_FIFO_out_0_port, cmd_valid_FIFO_out, cmd_ready_FIFO_out : std_logic;

begin
   
   Inst_PreProcessor : PreProcessor_2 port map( clk => clk, rst => rst, 
                           pdi_data(31) => pdi_data(31), pdi_data(30) => 
                           pdi_data(30), pdi_data(29) => pdi_data(29), 
                           pdi_data(28) => pdi_data(28), pdi_data(27) => 
                           pdi_data(27), pdi_data(26) => pdi_data(26), 
                           pdi_data(25) => pdi_data(25), pdi_data(24) => 
                           pdi_data(24), pdi_data(23) => pdi_data(23), 
                           pdi_data(22) => pdi_data(22), pdi_data(21) => 
                           pdi_data(21), pdi_data(20) => pdi_data(20), 
                           pdi_data(19) => pdi_data(19), pdi_data(18) => 
                           pdi_data(18), pdi_data(17) => pdi_data(17), 
                           pdi_data(16) => pdi_data(16), pdi_data(15) => 
                           pdi_data(15), pdi_data(14) => pdi_data(14), 
                           pdi_data(13) => pdi_data(13), pdi_data(12) => 
                           pdi_data(12), pdi_data(11) => pdi_data(11), 
                           pdi_data(10) => pdi_data(10), pdi_data(9) => 
                           pdi_data(9), pdi_data(8) => pdi_data(8), pdi_data(7)
                           => pdi_data(7), pdi_data(6) => pdi_data(6), 
                           pdi_data(5) => pdi_data(5), pdi_data(4) => 
                           pdi_data(4), pdi_data(3) => pdi_data(3), pdi_data(2)
                           => pdi_data(2), pdi_data(1) => pdi_data(1), 
                           pdi_data(0) => pdi_data(0), pdi_valid => pdi_valid, 
                           pdi_ready => pdi_ready, sdi_data(31) => sdi_data(31)
                           , sdi_data(30) => sdi_data(30), sdi_data(29) => 
                           sdi_data(29), sdi_data(28) => sdi_data(28), 
                           sdi_data(27) => sdi_data(27), sdi_data(26) => 
                           sdi_data(26), sdi_data(25) => sdi_data(25), 
                           sdi_data(24) => sdi_data(24), sdi_data(23) => 
                           sdi_data(23), sdi_data(22) => sdi_data(22), 
                           sdi_data(21) => sdi_data(21), sdi_data(20) => 
                           sdi_data(20), sdi_data(19) => sdi_data(19), 
                           sdi_data(18) => sdi_data(18), sdi_data(17) => 
                           sdi_data(17), sdi_data(16) => sdi_data(16), 
                           sdi_data(15) => sdi_data(15), sdi_data(14) => 
                           sdi_data(14), sdi_data(13) => sdi_data(13), 
                           sdi_data(12) => sdi_data(12), sdi_data(11) => 
                           sdi_data(11), sdi_data(10) => sdi_data(10), 
                           sdi_data(9) => sdi_data(9), sdi_data(8) => 
                           sdi_data(8), sdi_data(7) => sdi_data(7), sdi_data(6)
                           => sdi_data(6), sdi_data(5) => sdi_data(5), 
                           sdi_data(4) => sdi_data(4), sdi_data(3) => 
                           sdi_data(3), sdi_data(2) => sdi_data(2), sdi_data(1)
                           => sdi_data(1), sdi_data(0) => sdi_data(0), 
                           sdi_valid => sdi_valid, sdi_ready => sdi_ready, 
                           key(31) => key_cipher_in_31_port, key(30) => 
                           key_cipher_in_30_port, key(29) => 
                           key_cipher_in_29_port, key(28) => 
                           key_cipher_in_28_port, key(27) => 
                           key_cipher_in_27_port, key(26) => 
                           key_cipher_in_26_port, key(25) => 
                           key_cipher_in_25_port, key(24) => 
                           key_cipher_in_24_port, key(23) => 
                           key_cipher_in_23_port, key(22) => 
                           key_cipher_in_22_port, key(21) => 
                           key_cipher_in_21_port, key(20) => 
                           key_cipher_in_20_port, key(19) => 
                           key_cipher_in_19_port, key(18) => 
                           key_cipher_in_18_port, key(17) => 
                           key_cipher_in_17_port, key(16) => 
                           key_cipher_in_16_port, key(15) => 
                           key_cipher_in_15_port, key(14) => 
                           key_cipher_in_14_port, key(13) => 
                           key_cipher_in_13_port, key(12) => 
                           key_cipher_in_12_port, key(11) => 
                           key_cipher_in_11_port, key(10) => 
                           key_cipher_in_10_port, key(9) => 
                           key_cipher_in_9_port, key(8) => key_cipher_in_8_port
                           , key(7) => key_cipher_in_7_port, key(6) => 
                           key_cipher_in_6_port, key(5) => key_cipher_in_5_port
                           , key(4) => key_cipher_in_4_port, key(3) => 
                           key_cipher_in_3_port, key(2) => key_cipher_in_2_port
                           , key(1) => key_cipher_in_1_port, key(0) => 
                           key_cipher_in_0_port, key_valid => 
                           key_valid_cipher_in, key_ready => 
                           key_ready_cipher_in, bdi(31) => 
                           bdi_cipher_in_31_port, bdi(30) => 
                           bdi_cipher_in_30_port, bdi(29) => 
                           bdi_cipher_in_29_port, bdi(28) => 
                           bdi_cipher_in_28_port, bdi(27) => 
                           bdi_cipher_in_27_port, bdi(26) => 
                           bdi_cipher_in_26_port, bdi(25) => 
                           bdi_cipher_in_25_port, bdi(24) => 
                           bdi_cipher_in_24_port, bdi(23) => 
                           bdi_cipher_in_23_port, bdi(22) => 
                           bdi_cipher_in_22_port, bdi(21) => 
                           bdi_cipher_in_21_port, bdi(20) => 
                           bdi_cipher_in_20_port, bdi(19) => 
                           bdi_cipher_in_19_port, bdi(18) => 
                           bdi_cipher_in_18_port, bdi(17) => 
                           bdi_cipher_in_17_port, bdi(16) => 
                           bdi_cipher_in_16_port, bdi(15) => 
                           bdi_cipher_in_15_port, bdi(14) => 
                           bdi_cipher_in_14_port, bdi(13) => 
                           bdi_cipher_in_13_port, bdi(12) => 
                           bdi_cipher_in_12_port, bdi(11) => 
                           bdi_cipher_in_11_port, bdi(10) => 
                           bdi_cipher_in_10_port, bdi(9) => 
                           bdi_cipher_in_9_port, bdi(8) => bdi_cipher_in_8_port
                           , bdi(7) => bdi_cipher_in_7_port, bdi(6) => 
                           bdi_cipher_in_6_port, bdi(5) => bdi_cipher_in_5_port
                           , bdi(4) => bdi_cipher_in_4_port, bdi(3) => 
                           bdi_cipher_in_3_port, bdi(2) => bdi_cipher_in_2_port
                           , bdi(1) => bdi_cipher_in_1_port, bdi(0) => 
                           bdi_cipher_in_0_port, bdi_valid => 
                           bdi_valid_cipher_in, bdi_ready => 
                           bdi_ready_cipher_in, bdi_pad_loc(3) => 
                           bdi_pad_loc_cipher_in_3_port, bdi_pad_loc(2) => 
                           bdi_pad_loc_cipher_in_2_port, bdi_pad_loc(1) => 
                           bdi_pad_loc_cipher_in_1_port, bdi_pad_loc(0) => 
                           bdi_pad_loc_cipher_in_0_port, bdi_valid_bytes(3) => 
                           bdi_valid_bytes_cipher_in_3_port, bdi_valid_bytes(2)
                           => bdi_valid_bytes_cipher_in_2_port, 
                           bdi_valid_bytes(1) => 
                           bdi_valid_bytes_cipher_in_1_port, bdi_valid_bytes(0)
                           => bdi_valid_bytes_cipher_in_0_port, bdi_size(2) => 
                           bdi_size_cipher_in_2_port, bdi_size(1) => 
                           bdi_size_cipher_in_1_port, bdi_size(0) => 
                           bdi_size_cipher_in_0_port, bdi_eot => 
                           bdi_eot_cipher_in, bdi_eoi => bdi_eoi_cipher_in, 
                           bdi_type(3) => bdi_type_cipher_in_3_port, 
                           bdi_type(2) => bdi_type_cipher_in_2_port, 
                           bdi_type(1) => bdi_type_cipher_in_1_port, 
                           bdi_type(0) => bdi_type_cipher_in_0_port, decrypt =>
                           decrypt_cipher_in, hash => hash_cipher_in, 
                           key_update => key_update_cipher_in, cmd(31) => 
                           cmd_FIFO_in_31_port, cmd(30) => cmd_FIFO_in_30_port,
                           cmd(29) => cmd_FIFO_in_29_port, cmd(28) => 
                           cmd_FIFO_in_28_port, cmd(27) => cmd_FIFO_in_27_port,
                           cmd(26) => cmd_FIFO_in_26_port, cmd(25) => 
                           cmd_FIFO_in_25_port, cmd(24) => cmd_FIFO_in_24_port,
                           cmd(23) => cmd_FIFO_in_23_port, cmd(22) => 
                           cmd_FIFO_in_22_port, cmd(21) => cmd_FIFO_in_21_port,
                           cmd(20) => cmd_FIFO_in_20_port, cmd(19) => 
                           cmd_FIFO_in_19_port, cmd(18) => cmd_FIFO_in_18_port,
                           cmd(17) => cmd_FIFO_in_17_port, cmd(16) => 
                           cmd_FIFO_in_16_port, cmd(15) => cmd_FIFO_in_15_port,
                           cmd(14) => cmd_FIFO_in_14_port, cmd(13) => 
                           cmd_FIFO_in_13_port, cmd(12) => cmd_FIFO_in_12_port,
                           cmd(11) => cmd_FIFO_in_11_port, cmd(10) => 
                           cmd_FIFO_in_10_port, cmd(9) => cmd_FIFO_in_9_port, 
                           cmd(8) => cmd_FIFO_in_8_port, cmd(7) => 
                           cmd_FIFO_in_7_port, cmd(6) => cmd_FIFO_in_6_port, 
                           cmd(5) => cmd_FIFO_in_5_port, cmd(4) => 
                           cmd_FIFO_in_4_port, cmd(3) => cmd_FIFO_in_3_port, 
                           cmd(2) => cmd_FIFO_in_2_port, cmd(1) => 
                           cmd_FIFO_in_1_port, cmd(0) => cmd_FIFO_in_0_port, 
                           cmd_valid => cmd_valid_FIFO_in, cmd_ready => 
                           cmd_ready_FIFO_in);
   Inst_Cipher : CryptoCore_2 port map( clk => clk, rst => rst, key(31) => 
                           key_cipher_in_31_port, key(30) => 
                           key_cipher_in_30_port, key(29) => 
                           key_cipher_in_29_port, key(28) => 
                           key_cipher_in_28_port, key(27) => 
                           key_cipher_in_27_port, key(26) => 
                           key_cipher_in_26_port, key(25) => 
                           key_cipher_in_25_port, key(24) => 
                           key_cipher_in_24_port, key(23) => 
                           key_cipher_in_23_port, key(22) => 
                           key_cipher_in_22_port, key(21) => 
                           key_cipher_in_21_port, key(20) => 
                           key_cipher_in_20_port, key(19) => 
                           key_cipher_in_19_port, key(18) => 
                           key_cipher_in_18_port, key(17) => 
                           key_cipher_in_17_port, key(16) => 
                           key_cipher_in_16_port, key(15) => 
                           key_cipher_in_15_port, key(14) => 
                           key_cipher_in_14_port, key(13) => 
                           key_cipher_in_13_port, key(12) => 
                           key_cipher_in_12_port, key(11) => 
                           key_cipher_in_11_port, key(10) => 
                           key_cipher_in_10_port, key(9) => 
                           key_cipher_in_9_port, key(8) => key_cipher_in_8_port
                           , key(7) => key_cipher_in_7_port, key(6) => 
                           key_cipher_in_6_port, key(5) => key_cipher_in_5_port
                           , key(4) => key_cipher_in_4_port, key(3) => 
                           key_cipher_in_3_port, key(2) => key_cipher_in_2_port
                           , key(1) => key_cipher_in_1_port, key(0) => 
                           key_cipher_in_0_port, key_valid => 
                           key_valid_cipher_in, key_ready => 
                           key_ready_cipher_in, bdi(31) => 
                           bdi_cipher_in_31_port, bdi(30) => 
                           bdi_cipher_in_30_port, bdi(29) => 
                           bdi_cipher_in_29_port, bdi(28) => 
                           bdi_cipher_in_28_port, bdi(27) => 
                           bdi_cipher_in_27_port, bdi(26) => 
                           bdi_cipher_in_26_port, bdi(25) => 
                           bdi_cipher_in_25_port, bdi(24) => 
                           bdi_cipher_in_24_port, bdi(23) => 
                           bdi_cipher_in_23_port, bdi(22) => 
                           bdi_cipher_in_22_port, bdi(21) => 
                           bdi_cipher_in_21_port, bdi(20) => 
                           bdi_cipher_in_20_port, bdi(19) => 
                           bdi_cipher_in_19_port, bdi(18) => 
                           bdi_cipher_in_18_port, bdi(17) => 
                           bdi_cipher_in_17_port, bdi(16) => 
                           bdi_cipher_in_16_port, bdi(15) => 
                           bdi_cipher_in_15_port, bdi(14) => 
                           bdi_cipher_in_14_port, bdi(13) => 
                           bdi_cipher_in_13_port, bdi(12) => 
                           bdi_cipher_in_12_port, bdi(11) => 
                           bdi_cipher_in_11_port, bdi(10) => 
                           bdi_cipher_in_10_port, bdi(9) => 
                           bdi_cipher_in_9_port, bdi(8) => bdi_cipher_in_8_port
                           , bdi(7) => bdi_cipher_in_7_port, bdi(6) => 
                           bdi_cipher_in_6_port, bdi(5) => bdi_cipher_in_5_port
                           , bdi(4) => bdi_cipher_in_4_port, bdi(3) => 
                           bdi_cipher_in_3_port, bdi(2) => bdi_cipher_in_2_port
                           , bdi(1) => bdi_cipher_in_1_port, bdi(0) => 
                           bdi_cipher_in_0_port, bdi_valid => 
                           bdi_valid_cipher_in, bdi_ready => 
                           bdi_ready_cipher_in, bdi_pad_loc(3) => 
                           bdi_pad_loc_cipher_in_3_port, bdi_pad_loc(2) => 
                           bdi_pad_loc_cipher_in_2_port, bdi_pad_loc(1) => 
                           bdi_pad_loc_cipher_in_1_port, bdi_pad_loc(0) => 
                           bdi_pad_loc_cipher_in_0_port, bdi_valid_bytes(3) => 
                           bdi_valid_bytes_cipher_in_3_port, bdi_valid_bytes(2)
                           => bdi_valid_bytes_cipher_in_2_port, 
                           bdi_valid_bytes(1) => 
                           bdi_valid_bytes_cipher_in_1_port, bdi_valid_bytes(0)
                           => bdi_valid_bytes_cipher_in_0_port, bdi_size(2) => 
                           bdi_size_cipher_in_2_port, bdi_size(1) => 
                           bdi_size_cipher_in_1_port, bdi_size(0) => 
                           bdi_size_cipher_in_0_port, bdi_eot => 
                           bdi_eot_cipher_in, bdi_eoi => bdi_eoi_cipher_in, 
                           bdi_type(3) => bdi_type_cipher_in_3_port, 
                           bdi_type(2) => bdi_type_cipher_in_2_port, 
                           bdi_type(1) => bdi_type_cipher_in_1_port, 
                           bdi_type(0) => bdi_type_cipher_in_0_port, decrypt_in
                           => decrypt_cipher_in, key_update => 
                           key_update_cipher_in, hash_in => hash_cipher_in, 
                           bdo(31) => bdo_cipher_out_31_port, bdo(30) => 
                           bdo_cipher_out_30_port, bdo(29) => 
                           bdo_cipher_out_29_port, bdo(28) => 
                           bdo_cipher_out_28_port, bdo(27) => 
                           bdo_cipher_out_27_port, bdo(26) => 
                           bdo_cipher_out_26_port, bdo(25) => 
                           bdo_cipher_out_25_port, bdo(24) => 
                           bdo_cipher_out_24_port, bdo(23) => 
                           bdo_cipher_out_23_port, bdo(22) => 
                           bdo_cipher_out_22_port, bdo(21) => 
                           bdo_cipher_out_21_port, bdo(20) => 
                           bdo_cipher_out_20_port, bdo(19) => 
                           bdo_cipher_out_19_port, bdo(18) => 
                           bdo_cipher_out_18_port, bdo(17) => 
                           bdo_cipher_out_17_port, bdo(16) => 
                           bdo_cipher_out_16_port, bdo(15) => 
                           bdo_cipher_out_15_port, bdo(14) => 
                           bdo_cipher_out_14_port, bdo(13) => 
                           bdo_cipher_out_13_port, bdo(12) => 
                           bdo_cipher_out_12_port, bdo(11) => 
                           bdo_cipher_out_11_port, bdo(10) => 
                           bdo_cipher_out_10_port, bdo(9) => 
                           bdo_cipher_out_9_port, bdo(8) => 
                           bdo_cipher_out_8_port, bdo(7) => 
                           bdo_cipher_out_7_port, bdo(6) => 
                           bdo_cipher_out_6_port, bdo(5) => 
                           bdo_cipher_out_5_port, bdo(4) => 
                           bdo_cipher_out_4_port, bdo(3) => 
                           bdo_cipher_out_3_port, bdo(2) => 
                           bdo_cipher_out_2_port, bdo(1) => 
                           bdo_cipher_out_1_port, bdo(0) => 
                           bdo_cipher_out_0_port, bdo_valid => 
                           bdo_valid_cipher_out, bdo_ready => 
                           bdo_ready_cipher_out, bdo_type(3) => 
                           bdo_type_cipher_out_3_port, bdo_type(2) => 
                           bdo_type_cipher_out_2_port, bdo_type(1) => 
                           bdo_type_cipher_out_1_port, bdo_type(0) => 
                           bdo_type_cipher_out_0_port, bdo_valid_bytes(3) => 
                           bdo_valid_bytes_cipher_out_3_port, 
                           bdo_valid_bytes(2) => 
                           bdo_valid_bytes_cipher_out_2_port, 
                           bdo_valid_bytes(1) => 
                           bdo_valid_bytes_cipher_out_1_port, 
                           bdo_valid_bytes(0) => 
                           bdo_valid_bytes_cipher_out_0_port, end_of_block => 
                           end_of_block_cipher_out, msg_auth_valid => 
                           msg_auth_valid, msg_auth_ready => msg_auth_ready, 
                           msg_auth => msg_auth);
   Inst_PostProcessor : PostProcessor_2 port map( clk => clk, rst => rst, 
                           bdo(31) => bdo_cipher_out_31_port, bdo(30) => 
                           bdo_cipher_out_30_port, bdo(29) => 
                           bdo_cipher_out_29_port, bdo(28) => 
                           bdo_cipher_out_28_port, bdo(27) => 
                           bdo_cipher_out_27_port, bdo(26) => 
                           bdo_cipher_out_26_port, bdo(25) => 
                           bdo_cipher_out_25_port, bdo(24) => 
                           bdo_cipher_out_24_port, bdo(23) => 
                           bdo_cipher_out_23_port, bdo(22) => 
                           bdo_cipher_out_22_port, bdo(21) => 
                           bdo_cipher_out_21_port, bdo(20) => 
                           bdo_cipher_out_20_port, bdo(19) => 
                           bdo_cipher_out_19_port, bdo(18) => 
                           bdo_cipher_out_18_port, bdo(17) => 
                           bdo_cipher_out_17_port, bdo(16) => 
                           bdo_cipher_out_16_port, bdo(15) => 
                           bdo_cipher_out_15_port, bdo(14) => 
                           bdo_cipher_out_14_port, bdo(13) => 
                           bdo_cipher_out_13_port, bdo(12) => 
                           bdo_cipher_out_12_port, bdo(11) => 
                           bdo_cipher_out_11_port, bdo(10) => 
                           bdo_cipher_out_10_port, bdo(9) => 
                           bdo_cipher_out_9_port, bdo(8) => 
                           bdo_cipher_out_8_port, bdo(7) => 
                           bdo_cipher_out_7_port, bdo(6) => 
                           bdo_cipher_out_6_port, bdo(5) => 
                           bdo_cipher_out_5_port, bdo(4) => 
                           bdo_cipher_out_4_port, bdo(3) => 
                           bdo_cipher_out_3_port, bdo(2) => 
                           bdo_cipher_out_2_port, bdo(1) => 
                           bdo_cipher_out_1_port, bdo(0) => 
                           bdo_cipher_out_0_port, bdo_valid => 
                           bdo_valid_cipher_out, bdo_ready => 
                           bdo_ready_cipher_out, end_of_block => 
                           end_of_block_cipher_out, bdo_type(3) => 
                           bdo_type_cipher_out_3_port, bdo_type(2) => 
                           bdo_type_cipher_out_2_port, bdo_type(1) => 
                           bdo_type_cipher_out_1_port, bdo_type(0) => 
                           bdo_type_cipher_out_0_port, bdo_valid_bytes(3) => 
                           bdo_valid_bytes_cipher_out_3_port, 
                           bdo_valid_bytes(2) => 
                           bdo_valid_bytes_cipher_out_2_port, 
                           bdo_valid_bytes(1) => 
                           bdo_valid_bytes_cipher_out_1_port, 
                           bdo_valid_bytes(0) => 
                           bdo_valid_bytes_cipher_out_0_port, msg_auth => 
                           msg_auth, msg_auth_ready => msg_auth_ready, 
                           msg_auth_valid => msg_auth_valid, cmd(31) => 
                           cmd_FIFO_out_31_port, cmd(30) => 
                           cmd_FIFO_out_30_port, cmd(29) => 
                           cmd_FIFO_out_29_port, cmd(28) => 
                           cmd_FIFO_out_28_port, cmd(27) => 
                           cmd_FIFO_out_27_port, cmd(26) => 
                           cmd_FIFO_out_26_port, cmd(25) => 
                           cmd_FIFO_out_25_port, cmd(24) => 
                           cmd_FIFO_out_24_port, cmd(23) => 
                           cmd_FIFO_out_23_port, cmd(22) => 
                           cmd_FIFO_out_22_port, cmd(21) => 
                           cmd_FIFO_out_21_port, cmd(20) => 
                           cmd_FIFO_out_20_port, cmd(19) => 
                           cmd_FIFO_out_19_port, cmd(18) => 
                           cmd_FIFO_out_18_port, cmd(17) => 
                           cmd_FIFO_out_17_port, cmd(16) => 
                           cmd_FIFO_out_16_port, cmd(15) => 
                           cmd_FIFO_out_15_port, cmd(14) => 
                           cmd_FIFO_out_14_port, cmd(13) => 
                           cmd_FIFO_out_13_port, cmd(12) => 
                           cmd_FIFO_out_12_port, cmd(11) => 
                           cmd_FIFO_out_11_port, cmd(10) => 
                           cmd_FIFO_out_10_port, cmd(9) => cmd_FIFO_out_9_port,
                           cmd(8) => cmd_FIFO_out_8_port, cmd(7) => 
                           cmd_FIFO_out_7_port, cmd(6) => cmd_FIFO_out_6_port, 
                           cmd(5) => cmd_FIFO_out_5_port, cmd(4) => 
                           cmd_FIFO_out_4_port, cmd(3) => cmd_FIFO_out_3_port, 
                           cmd(2) => cmd_FIFO_out_2_port, cmd(1) => 
                           cmd_FIFO_out_1_port, cmd(0) => cmd_FIFO_out_0_port, 
                           cmd_valid => cmd_valid_FIFO_out, cmd_ready => 
                           cmd_ready_FIFO_out, do_data(31) => do_data(31), 
                           do_data(30) => do_data(30), do_data(29) => 
                           do_data(29), do_data(28) => do_data(28), do_data(27)
                           => do_data(27), do_data(26) => do_data(26), 
                           do_data(25) => do_data(25), do_data(24) => 
                           do_data(24), do_data(23) => do_data(23), do_data(22)
                           => do_data(22), do_data(21) => do_data(21), 
                           do_data(20) => do_data(20), do_data(19) => 
                           do_data(19), do_data(18) => do_data(18), do_data(17)
                           => do_data(17), do_data(16) => do_data(16), 
                           do_data(15) => do_data(15), do_data(14) => 
                           do_data(14), do_data(13) => do_data(13), do_data(12)
                           => do_data(12), do_data(11) => do_data(11), 
                           do_data(10) => do_data(10), do_data(9) => do_data(9)
                           , do_data(8) => do_data(8), do_data(7) => do_data(7)
                           , do_data(6) => do_data(6), do_data(5) => do_data(5)
                           , do_data(4) => do_data(4), do_data(3) => do_data(3)
                           , do_data(2) => do_data(2), do_data(1) => do_data(1)
                           , do_data(0) => do_data(0), do_valid => do_valid, 
                           do_last => do_last, do_ready => do_ready);
   Inst_Header_Fifo : fwft_fifo_G_W32_G_LOG2DEPTH2 port map( clk => clk, rst =>
                           rst, din(31) => cmd_FIFO_in_31_port, din(30) => 
                           cmd_FIFO_in_30_port, din(29) => cmd_FIFO_in_29_port,
                           din(28) => cmd_FIFO_in_28_port, din(27) => 
                           cmd_FIFO_in_27_port, din(26) => cmd_FIFO_in_26_port,
                           din(25) => cmd_FIFO_in_25_port, din(24) => 
                           cmd_FIFO_in_24_port, din(23) => cmd_FIFO_in_23_port,
                           din(22) => cmd_FIFO_in_22_port, din(21) => 
                           cmd_FIFO_in_21_port, din(20) => cmd_FIFO_in_20_port,
                           din(19) => cmd_FIFO_in_19_port, din(18) => 
                           cmd_FIFO_in_18_port, din(17) => cmd_FIFO_in_17_port,
                           din(16) => cmd_FIFO_in_16_port, din(15) => 
                           cmd_FIFO_in_15_port, din(14) => cmd_FIFO_in_14_port,
                           din(13) => cmd_FIFO_in_13_port, din(12) => 
                           cmd_FIFO_in_12_port, din(11) => cmd_FIFO_in_11_port,
                           din(10) => cmd_FIFO_in_10_port, din(9) => 
                           cmd_FIFO_in_9_port, din(8) => cmd_FIFO_in_8_port, 
                           din(7) => cmd_FIFO_in_7_port, din(6) => 
                           cmd_FIFO_in_6_port, din(5) => cmd_FIFO_in_5_port, 
                           din(4) => cmd_FIFO_in_4_port, din(3) => 
                           cmd_FIFO_in_3_port, din(2) => cmd_FIFO_in_2_port, 
                           din(1) => cmd_FIFO_in_1_port, din(0) => 
                           cmd_FIFO_in_0_port, din_valid => cmd_valid_FIFO_in, 
                           din_ready => cmd_ready_FIFO_in, dout(31) => 
                           cmd_FIFO_out_31_port, dout(30) => 
                           cmd_FIFO_out_30_port, dout(29) => 
                           cmd_FIFO_out_29_port, dout(28) => 
                           cmd_FIFO_out_28_port, dout(27) => 
                           cmd_FIFO_out_27_port, dout(26) => 
                           cmd_FIFO_out_26_port, dout(25) => 
                           cmd_FIFO_out_25_port, dout(24) => 
                           cmd_FIFO_out_24_port, dout(23) => 
                           cmd_FIFO_out_23_port, dout(22) => 
                           cmd_FIFO_out_22_port, dout(21) => 
                           cmd_FIFO_out_21_port, dout(20) => 
                           cmd_FIFO_out_20_port, dout(19) => 
                           cmd_FIFO_out_19_port, dout(18) => 
                           cmd_FIFO_out_18_port, dout(17) => 
                           cmd_FIFO_out_17_port, dout(16) => 
                           cmd_FIFO_out_16_port, dout(15) => 
                           cmd_FIFO_out_15_port, dout(14) => 
                           cmd_FIFO_out_14_port, dout(13) => 
                           cmd_FIFO_out_13_port, dout(12) => 
                           cmd_FIFO_out_12_port, dout(11) => 
                           cmd_FIFO_out_11_port, dout(10) => 
                           cmd_FIFO_out_10_port, dout(9) => cmd_FIFO_out_9_port
                           , dout(8) => cmd_FIFO_out_8_port, dout(7) => 
                           cmd_FIFO_out_7_port, dout(6) => cmd_FIFO_out_6_port,
                           dout(5) => cmd_FIFO_out_5_port, dout(4) => 
                           cmd_FIFO_out_4_port, dout(3) => cmd_FIFO_out_3_port,
                           dout(2) => cmd_FIFO_out_2_port, dout(1) => 
                           cmd_FIFO_out_1_port, dout(0) => cmd_FIFO_out_0_port,
                           dout_valid => cmd_valid_FIFO_out, dout_ready => 
                           cmd_ready_FIFO_out);

end SYN_structure;

library IEEE;

use IEEE.std_logic_1164.all;
entity SELECT_OP is
   generic ( num_inputs, input_width : integer );
   port(
      DATA : in std_logic_vector( num_inputs  * input_width - 1 downto 0 );
      CONTROL : in std_logic_vector( num_inputs - 1 downto 0 );
      Z : out std_logic_vector( input_width - 1 downto 0 )
   );
end SELECT_OP;

architecture RTL of SELECT_OP is
begin

   process ( DATA, CONTROL )
      variable index, high, low : integer;
   begin
   
      --  Initialize variables
      index := 0;
      
      -- Loop over the values of the control inputs
      for_loop : for i in CONTROL'range loop
      
         if ( CONTROL(i) = '1' ) then
         
            index := i;
            exit for_loop;
            
         end if;
         
      end loop;
      
      -- Store the corresponding data lines into the output
      low := input_width * index;
      high := low + input_width - 1;
      Z <= DATA( high downto low );
   
   end process;
   
end RTL;

library IEEE;

use IEEE.std_logic_1164.all;

entity SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT is
   generic ( ac_as_q, ac_as_qn, sc_ss_q : integer );
   port(
      clear, preset, enable, data_in, synch_clear, synch_preset, synch_toggle, 
         synch_enable, next_state, clocked_on : in std_logic;
      Q, QN : buffer std_logic
   );
end SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT;

architecture RTL of SYNOPSYS_BASIC_SEQUENTIAL_ELEMENT is
begin

   process ( preset, clear, enable, data_in, clocked_on )
   begin
   
            -- Check the value of inputs (asynchronous first)
            if ( ( ( preset /= '1' ) and ( preset /= '0' ) ) or ( ( clear /= 
                     '1' ) and ( clear /= '0' ) )  ) then
               Q <= 'X';
            elsif ( clear = '1' and preset = '1' ) then
               case ac_as_q is
                  when 2 =>
                     Q <= '1';
                  when 1 =>
                     Q <= '0';
                  when others =>
                     Q <= 'X';
               end case;
               case ac_as_qn is
                  when 2 =>
                     QN <= '1';
                  when 1 =>
                     QN <= '0';
                  when others =>
                     QN <= 'X';
               end case;
            elsif ( clear = '1' ) then
               Q <= '0';
            elsif ( preset = '1' ) then
               Q <= '1';
            elsif ( ( enable /= '1' ) and ( enable /= '0' ) ) then
               Q <= 'X';
            elsif ( enable = '1' ) then
               Q <= data_in;
            elsif ( ( clocked_on /= '1' ) and ( clocked_on /= '0' ) ) then
               Q <= 'X';
            elsif ( clocked_on'event and clocked_on = '1' ) then
         if ( ( ( synch_preset /= '1' ) and ( synch_preset /= '0' ) ) or ( ( 
                  synch_clear /= '1' ) and ( synch_clear /= '0' ) )  ) then
            Q <= 'X';
         elsif ( synch_clear = '1' and synch_preset = '1' ) then
            case sc_ss_q is
               when 2 =>
                  Q <= '1';
               when 1 =>
                  Q <= '0';
               when others =>
                  Q <= 'X';
            end case;
         elsif ( synch_clear = '1' ) then
            Q <= '0';
         elsif ( synch_preset = '1' ) then
            Q <= '1';
         elsif ( ( ( synch_toggle /= '1' ) and ( synch_toggle /= '0' ) ) or ( (
                  synch_enable /= '1' ) and ( synch_enable /= '0' ) )  ) then
            Q <= 'X';
         elsif ( synch_enable = '1' and synch_toggle = '1' ) then
            Q <= 'X';
         elsif ( synch_toggle = '1' ) then
            Q <= QN;
         elsif ( synch_enable = '1' ) then
            Q <= next_state;
         end if;
      end if;
   
   end process;

end RTL;
